���      �xgboost.sklearn��XGBClassifier���)��}�(�use_label_encoder�N�n_estimators�Kd�	objective��multi:softprob��	max_depth�N�
max_leaves�N�max_bin�N�grow_policy�N�learning_rate�N�	verbosity�N�booster�N�tree_method�N�gamma�N�min_child_weight�N�max_delta_step�N�	subsample�N�sampling_method�N�colsample_bytree�N�colsample_bylevel�N�colsample_bynode�N�	reg_alpha�N�
reg_lambda�N�scale_pos_weight�N�
base_score�N�missing�G�      �num_parallel_tree�N�random_state�N�n_jobs�N�monotone_constraints�N�interaction_constraints�N�importance_type�N�gpu_id�N�validate_parameters�N�	predictor�N�enable_categorical���feature_types�N�max_cat_to_onehot�N�max_cat_threshold�N�eval_metric�N�early_stopping_rounds�N�	callbacks�N�classes_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h2�dtype����i4�����R�(K�<�NNNJ����J����K t�b�C          �t�b�
n_classes_�K�_Booster��xgboost.core��Booster���)��}�(�handle��builtins��	bytearray���B@ {L       Config{L       learner{L       generic_param{L       fail_on_invalid_gpu_idSL       0L       gpu_idSL       -1L       n_jobsSL       0L       nthreadSL       0L       random_stateSL       0L       seedSL       0L       seed_per_iterationSL       0L       validate_parametersSL       1}L       gradient_booster{L       gbtree_model_param{L       num_parallel_treeSL       1L       	num_treesSL       300L       size_leaf_vectorSL       0}L       gbtree_train_param{L       	predictorSL       autoL       process_typeSL       defaultL       tree_methodSL       exactL       updaterSL       grow_colmaker,pruneL       updater_seqSL       grow_colmaker,prune}L       nameSL       gbtreeL       specified_updaterFL       updater{L       grow_colmaker{L       colmaker_train_param{L       default_directionSL       learnL       opt_dense_colSL       1}L       train_param{L       alphaSL       0L       	cache_optSL       1L       colsample_bylevelSL       1L       colsample_bynodeSL       1L       colsample_bytreeSL       1L       etaSL       0.300000012L       gammaSL       0L       grow_policySL       	depthwiseL       interaction_constraintsSL        L       lambdaSL       1L       learning_rateSL       0.300000012L       max_binSL       256L       max_cat_thresholdSL       64L       max_cat_to_onehotSL       4L       max_delta_stepSL       0L       	max_depthSL       6L       
max_leavesSL       0L       min_child_weightSL       1L       min_split_lossSL       0L       monotone_constraintsSL       ()L       refresh_leafSL       1L       	reg_alphaSL       0L       
reg_lambdaSL       1L       sampling_methodSL       uniformL       sketch_ratioSL       2L       sparse_thresholdSL       0.20000000000000001L       	subsampleSL       1}}L       prune{L       train_param{L       alphaSL       0L       	cache_optSL       1L       colsample_bylevelSL       1L       colsample_bynodeSL       1L       colsample_bytreeSL       1L       etaSL       0.300000012L       gammaSL       0L       grow_policySL       	depthwiseL       interaction_constraintsSL        L       lambdaSL       1L       learning_rateSL       0.300000012L       max_binSL       256L       max_cat_thresholdSL       64L       max_cat_to_onehotSL       4L       max_delta_stepSL       0L       	max_depthSL       6L       
max_leavesSL       0L       min_child_weightSL       1L       min_split_lossSL       0L       monotone_constraintsSL       ()L       refresh_leafSL       1L       	reg_alphaSL       0L       
reg_lambdaSL       1L       sampling_methodSL       uniformL       sketch_ratioSL       2L       sparse_thresholdSL       0.20000000000000001L       	subsampleSL       1}}}}L       learner_model_param{L       
base_scoreSL       5E-1L       boost_from_averageSL       1L       	num_classSL       3L       num_featureSL       8L       
num_targetSL       1}L       learner_train_param{L       boosterSL       gbtreeL       disable_default_eval_metricSL       0L       dsplitSL       autoL       	objectiveSL       multi:softprob}L       metrics[#L       {L       nameSL       mlogloss}L       	objective{L       nameSL       multi:softprobL       softmax_multiclass_param{L       	num_classSL       3}}}L       version[#L       iii}L       Model{L       learner{L       
attributes{L       best_iterationSL       99L       best_ntree_limitSL       100}L       feature_names[#L       SL       BALANCESL       	PURCHASESSL       PURCHASES_FREQUENCYSL       CASH_ADVANCE_FREQUENCYSL       CASH_ADVANCE_TRXSL       PURCHASES_TRXSL       PAYMENTSSL       MINIMUM_PAYMENTSL       feature_types[#L       SL       floatSL       floatSL       floatSL       floatSL       floatSL       floatSL       floatSL       floatL       gradient_booster{L       model{L       gbtree_model_param{L       num_parallel_treeSL       1L       	num_treesSL       300L       size_leaf_vectorSL       0}L       	tree_info[#L      ,i iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iii iiL       trees[#L      ,{L       base_weights[$d#L       _��"=?��Ӿ�f�>�O�?��9�Af>�n�,C?�B?|-�?�l�2���ip�?�M��g,���=?�i�?#�~?���>�1�?�;?�
�?��ÿ:�z�Ŗ�?d.+�N!?��\���P�Z�ۿ5>��>�����?Ri4?dS==ǳ��?�
��=�(�蒉>��׿7g+?�tQ>͛5>�3�*�?���?���*��>L�˾���>�(�zƋ�8�ɿ4�`�(T5�IqZ?dS>�ڈ?�ډ����?[m�>�m���m�?��)?�ֿ)�̿?$�?���*T(���?:.��9����m�?-kZ?��"<k-%?T'�?[m��Q�d��k��5�b?��?�@�?�Wӽ�\e?[m�����/^����#?6T���m��L>�m�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       _                                                L       idi L       left_children[$l#L       _               	                                 ����   !����   #����   %����   '   )   +   -   /   1   3   5   7   9����   ;����   =   ?   A   C   E   G   I   K   M   O   Q   S   U����   W   Y   [   ]��������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       _D��&B��pC��#A�@@4� B�� C���@�e?��p@��(?� A�b`C ,B��A��"@��4    ?�L�    ?�^�    @��    @�ʀBG,A�_|Ao5�AC��@�A�:Y?0��@ĺ@
o�    ?��    @
�?[m�? >v  At,�Al<�?1N�@`@߯t@�H�@�5�A�AE    ?��AUQA��?��"                                                                                                                                                                    L       parents[$l#L       _���                                                           	   	   
   
                                                                                                                 "   "   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   2   2   3   3   4   4   5   5L       right_children[$l#L       _               
                                  ����   "����   $����   &����   (   *   ,   .   0   2   4   6   8   :����   <����   >   @   B   D   F   H   J   L   N   P   R   T   V����   X   Z   \   ^��������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       _��fT�[Q�>��.;�l�D�8>ג�=Ox�?|� >��6���$� �*�JA��n?v�?����[&>�儿nwI>�M�T��>ԭL�,�>�?�(��f��d���2�>�?�@?��侑?��V�^��&�t��V��>�������Jm����������о�T�@JE�?)�&?��j><��+���BPh���L��?���0�H?2V�>�<��]�X�Y1A�I���q�9>���=��
>�����>��:>�:��<>�B�>�F5�K���e_�>8Q�Ld���>_k�^�E��;>Pm>�n);�>~��>��;�{ݬ����ZH�>_�>�M�>��ʽ=>��:���L�Rq���8�>Z���<�.[U>�:L       split_indices[$l#L       _                                                                                                                                                                                                                                                                                                                                                        L       
split_type[$U#L       _                                                                                               L       sum_hessian[$d#L       _E[q�DLq�E(UUBgqD=��E��DUUB
��A��A���D8��Dݎ8C��Cw��C���B�@8�A8�Ac�8AUUA?��B�q�D"qD�*�C#qB�8�C�8�Ck��A?��CqC8�A�q�A8�?�8@�8@Gq@�q@*��B�qD���B��8BQ�B�UTBWqB%UUAÎ8C���CS��A���@���@��B��Bx�@�8�C�A��8@�8@��@Gq@c�8@c�8@�q�?���?���?���B
��BS�8B�qD��A*��B\q�A��8A���Bڪ�?���AUUB1�A��A��@��A�qA�8�Cv8�A\q�CF8�Ac�8Aq�?���@*��B%UUBN8�B5UUA�q@Gq?���L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       95L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       I��"=�7�?.���8�?[m�>��m?��"�?�Fs���?"'�>���?��|�0t9>+*ȿ@�?-kZ����?oh��;6�?���?�_�?�׹�;4"�f�=���>��/�1Q���>5���?�y��;�?+>���?����q?M�>�m�?���?�?��y�<�x��m�?&ֿ�;��m��(T+���?�5�5Y����P�4P%>��ڿM�>�m�>�Ƈ?� Y�#����*��Es?B��i��?G�?S��?���+ܾ,����?�  =���?gSG?C}�?�eL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       I                                     L       idiL       left_children[$l#L       I            ����   	   ����                                 !   #   %   '����   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C��������   E   G��������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       ID�'EAP/ C���@�s     Ck��Br��    A��B{vC!� A�a\A>Q @=� @�l�A��`BU�B%�A�Aa,=6� Ac�`    ?83 @��>�{�@�5O?NP A�1�?�b�?��A-�^A$��A�olA���?���@�        @���@jV                                                                                                                                 L       parents[$l#L       I���                                               	   	   
   
                                                                                                                                   !   !   "   "   #   #   $   $   '   '   (   (L       right_children[$l#L       I            ����   
   ����                                  "   $   &   (����   *   ,   .   0   2   4   6   8   :   <   >   @   B   D��������   F   H��������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       I���1?Հ�?oh<��P>��;��I�`�e;��Z??��<ޜb>�=�>�H�>Ĺ�����>���o��?O&ԿK�t?���?7�޿/��>�6@��?�.��
>�q�����x%��g���h��[�:���+?K�^>���.�f�$��>�:>��Ⱦ�/�>����b�*��;>GCξ���;�I���8Q�>1s�Y�ͽ�NǾX`-=��l�1��>�:>w>��C�㼬v�����>i�ڽ�P>ox�>~[\>�zN�MT��O�t�>���<��l>�ˑ>j��>�yQL       split_indices[$l#L       I                                                                                                                                                                                                                                                                        L       
split_type[$U#L       I                                                                         L       sum_hessian[$d#L       IE[q�D�8�DપDժ�@�8�D��D0UUD�qCDq�C�q�D4�Ba�D"8�C�8B�8C�qBJ��CQ�D UUBq�A���CW�8Cت�C�A\q�AqA�8C]UTB��A��8B�CUUB��B��C�q�AꪪAq�?���A��B(�C-UUCq�?���@GqA*��?���@�8@��AÎ8CQUUA?��BUUBn8�Aq�?���@�8�A�8�B���B_��A�UUBGqA��B%UUC�UUC68�A��8A8�?�8@���Ax�A�UTA���C��L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       73L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       q9F�@?��/��u^?�B5�W�B=�ڿ\�?�F㾄�;?/���p�?1���X>��/�#�/?�$I�b��>/�����?x��ڊ���=�څ?n�������o��~^�?+���4�N?��,?u�>?Vd���L>�NľzƋ�`0>�ܰ?�Y>�qO��ֿ%����?��?�#�<� �?����8>��r�����i��4D>���,��?�p��C'����*�����^�8?��x?�ڦ?�@~�i�?����m������W?<`���m�>u���L�Ͽ3c
>u?�k[?;Q+�Sܳ?u����m��.d����P?����%D>�˖?�k[�Sܳ����2�>�}g��i��.��06>�m���_@���5͠���?,h}?�ƽ�>�m�����ƽ~ؓ�>iʿ#ʿ4��>~=�>jc�+h<L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       q                                                         L       idiL       left_children[$l#L       q               	                                    !   #   %   '����   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I����   K   M   O   Q��������   S   U   W   Y   [   ]   _   a   c����   e   g   i   k   m   o����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       qD��B��0C�z�B�:�A�JC}h�A�@B9�@@J5HA2�?��hB�<B�Q�Ax�A]s@A>�@�K�?��R@)��@ ��    ?�L�?��MB�L�A�VB�X�A��@���ATAV<�@CZ ?�� @�p(@v�?��@
�?l�?�x    ?�� ?Î$@�A�?�p        A���A���@�H�@a�XB5��@��pAd ?�v�@�<    @@�P?�CA�#Z?��@A�=?#t                                                                                                                                                                                                                 L       parents[$l#L       q���                                                           	   	   
   
                                                                                                                                   !   !   "   "   #   #   $   $   %   %   '   '   (   (   )   )   *   *   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   7   7   8   8   9   9   :   :   ;   ;   <   <L       right_children[$l#L       q               
                                     "   $   &   (����   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J����   L   N   P   R��������   T   V   X   Z   \   ^   `   b   d����   f   h   j   l   n   p����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       q�[��?���.$�;�l�=��p��Q��Kv�?N��>��6@5#Z�] �?��>� |�;�>����� g�o��>�8���E��0&@�3�?�����	>�[Y�o��>�(�>�]f���$?v�=����'��>Ыq?��@ >�?��r?�0�`�5�m=�<�{8F��v/�c�ݿ p�t�>8Q뿏��]��=TT�>U�?��P?�g>�����'�T���O�?O��>�"�����Ұݾݑ��QB>���>��.>�1��>���<�-zU�0	6>b���<=�t��'�K�u�WC�=�t�>�n>`�ν~<>�t��<��;�QE���N�>�Fy�FQ�>	��>�n�~<�󺣾V�,>���7��k�St>�:���'�K�Z)���C�>N��>����t�>�:�<�>�T���Y�d~�+Č�X��=�q�d��M�IL       split_indices[$l#L       q                                                                                                                                                                                                                                                                                                                                                                                                                     L       
split_type[$U#L       q                                                                                                                 L       sum_hessian[$d#L       qE[q�D18�E/#�D#8�B_��D��8D���Dq�A��A��8B8�C�UUDmq�BqD���D��A��A*��A��8A�q@c�8A���@c�8C��B��DqCª�A��8A���C���Ds��D
�8B1�@��A���@�q@�8�A��@8�A1�@��@�qA�8�?�8?�8C��8B�UUA8�B���C���C8q�B�8C��@��A8�Ax�@��C[��CS��BO��Df��D��A��B(�@8�@�8�?���AqA8�@�q�?���?�8@*��@��Ac�8?�8AUU@c�8@8�?�8@�8�?���AÎ8A?��C{qAʪ�B%UUAUU@8�AGqBS�8C�UUBª�B���B��A*��B�8�@*��C�q�@Gq@�8�A\q�?�8?���@�8�BÎ8B�q�B���B���B�A\q�D8�C��8L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       113L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       o�]��?C���߱_�7�?h���
�>�1��P�?ND3>���?��& s��u�?CJ;��@`��W�(��>}*?X�l?j����A�?i>?�H�'�1��ա>��n�H7?i��=�K뽏��%��l�R?	E���ֿ+o�?:^���^\?f_�>����?qԱ��J?T�:?4�U?f?�j�>ѐ��(��>Z�?v�	�?�Z���9=�z��!ts?nMt��]���6?Yھ���>�&��(=��İ���>�
>L�?bf\��c=��?(��?|A��}�?c��>����ڿ�?T�^?�w���?[�C?v�����?H�_����?���>d!�)Ǒ���?#X!�x[<����r�>w�P?y
�>�Hu��Ha��|?�M�'>����>�w�?yvi?>�Z��gH?MQJ��E��#�׽:�U?����=ɬ5��|�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       o                                                        L       idiL       left_children[$l#L       o               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C������������   E   G   I   K   M   O   Q   S��������   U   W����   Y   [   ]   _   a   c����   e   g   i   k����   m������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       oD���C��C>�BGb{B#�A�` B��ZA2D�?F� B#��=  @�� BG��A�e\A�(@���;Ԁ ?��?G� @(6@A�#?�� =N@ @G @�p�A#0�A7��@}� @��Ao=�=� @��?Ġ�>�Y>            =�� @1:~?:r�>x� @��@~��@\�p?         ?� @�/�    >��@�K�@�6@�-�@c�@d.�    @V�@E�A ͆A�    >���                                                                                                                                                                                                L       parents[$l#L       o���                                                           	   	   
   
                                                                                                                                         !   !   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   /   /   0   0   2   2   3   3   4   4   5   5   6   6   7   7   9   9   :   :   ;   ;   <   <   >   >L       right_children[$l#L       o               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D������������   F   H   J   L   N   P   R   T��������   V   X����   Z   \   ^   `   b   d����   f   h   j   l����   n������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       o�P7�Gh>��.���$� �*>�dL>fw�W���o�x�Sԭ���
?O����>�]�??�Ⱦ�[&��l��pR��O�y�,�>Fz:>~|��F@9��`g=�X��2�?m�8?��h?���@F�t�����&�nr�M�%>_�Ӿkѿj�Ⱦ��!�Jm�R T?PH�?gyg�F��^͘>�L�=�zc?�#S�5 >��߾�.�?����<�`<��?O��?)S��Ҿ��,?7��<2+>�R�I��?P#��!��=�z�=5�r>���!��<���>JN�>�ZC�KU>���=ۖ��?�>">�)��\>���>�꽷�d>p�?����>���=����K�H��u>D[�']:;��߾;�=���>�l�=�V�^����B>�*I�H�����Y=�)>��s>d�����>va��� T�D�ϼ` >,Ѣ����<�ھ�]L       split_indices[$l#L       o                                                                                                                                                                                                                                                                                                                                                                                                                L       
split_type[$U#L       o                                                                                                               L       sum_hessian[$d#L       oEQ@�D���E�FC%�RD�!SDӰ#C��B�{pB%�fC7S�DVm�D��C�p�C;�dC�tB&o}B�C�@V�RB��Bɕ�B�B�� D6��D�A�Ai2B�yCq��C�DB�C�B��,A�wvA4�
@��B��1?�?���B�@�)�@/XB��BkJ�A���B"�B���D6�?�i�D�b�Aoh3@���A(Z)Bd��A�z�A͟�CW��C�j?��(A�- A~��B�/OB}��B�?�@tF=A�\0A26�@Ѧ	@��
@^s�?���A2�A��?��@�??��?�BF��BAs�B]q�@]�qA��@'�B1@-�RB��Y?���D�qEA�_@��rA*�z?��nA�A��7A���@p�Ad��A�MZ@R��COA�A.#FC5?�+A�jNAP�,@6�DB*�mB?�2B,$vA��j?���@*|L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       111L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       Q:9��#�p? �!�$��?-����?�?��+7����>��?d-��=� C>�˱?jEͿ=ԥL�'��G4���Cb>��~�_?�?C�?}d��'���P����>�?��)�l�����>�I�?Ґ� O�>�?����"?��=A�^?.��>��T?_��?�I?~�d�)��=ԫ��m�?0�ӿR <ĞH����>��׿+km�p�D�����μ���z?"U�� 9����� ��?D!�>�ԗ?����Ի?
�V>F�?X˾���>���>�N?aJ�<�_�? ��?W�?z>�%c*?-��?�?�TL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       Q                                         L       idiL       left_children[$l#L       Q               	      ����   ��������                           !   #   %   '   )   +   -   /   1   3   5����   7   9����   ;   =   ?   A   C   E   G   I   K   M   O������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       QD��WA��CY��@�� >� A:��B��    Aw6,        @��@@��B��T@�� @�0@���>�[ @�$h@4@&@g��B�wB 9XA;�@?v� ?)��@JB_>�P�@�>�\�    >��P?�4y    ?��@
ʸ=ԇ A,@���AVoA��P@���@�� ?��2>�`                                                                                                                                                 L       parents[$l#L       Q���                                                                                                                                                                                     "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,L       right_children[$l#L       Q               
      ����   ��������                            "   $   &   (   *   ,   .   0   2   4   6����   8   :����   <   >   @   B   D   F   H   J   L   N   P������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       Q���1?Հ���n<��P?���?N��?&l��MuI�Z=�L�>��]>�ΐ���?->��>Ĺ����@0}�>.R?ax>?��>���J�K�ǮO@��?-��?kE�>�ŵ@.ν+]�?���v>4�����t@G�?|�l?�,=󦔽^<&�#?���>����ʡa�gʆ�K��<02g��>T��?/4;��$�ħ>v�M���^��1S��|� O�>B�I�@Di��S�@��>k[�=��>����$2z>&y4=0�Y>�����=�=�Q$>wb>�,�;�r�>A%�>6��>�%F�Fw >P�c>.�$>���L       split_indices[$l#L       Q                                                                                                                                                                                                                                                                                                   L       
split_type[$U#L       Q                                                                                 L       sum_hessian[$d#L       QERZDD�  D�gD�fO@�ѣCPفDљ7D�=�C1B�@��@�MC�
BE!�Dc>�D?�Cj�B`�C��A���A�i�A��1CY�eD,ׄC���C�@B��AV3@��A�;C�@c�Ax�!A��?��A�)VA���@�X�C&�gBK��B璉D�BW��CK��@���C�j�B��Q?�$?A2-�@@��h?�w@��pA�TC��@/��AY2�?�2�?�Ҟ@�D�Al�Au�Aj�H@S
j?��@�C�X@���A�߂AԸiBQ�B�%�C�1C��2A�zA�'|Bd/C��?�'�@��@�w�C�<�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       81L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       q;�?9T澕�m?YBF���QKw�1N?g�����>��H� �>��o�q�����ҿ8�?tnm=�(��\k?߷?(���7��"���?"�ھ���e*�
8޾9U���a��x�&��?�?z��??@̾<�h>N�ݾ��o?]�� F�?6�?���]�rI>/ξ�7�?h޽� ~�5�?E����?
�F��S>z��7���� ��>FO־׃�� �v<�\ݿ&ޮ��Z�?9�H<��?���?9Z�=i�?eȖ>�����=�?�s�햢�X���#�>�4�?|��?��v>�wt���=cy���6?4z����=51j���4~C��N�?W=R�#�5<�a?Cz>���>@Ɖ�
�?:v���>3�r�:�>���5=9z]�#q��Ύ?T�e���5п"_:=<�i?w�?��u�*)u?
�ֿ�wL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       q                                                         L       idiL       left_children[$l#L       q               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;����   =   ?   A   C   E   G   I����   K����   M   O   Q��������   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       qD3�B�"�C0�B7ppA�{2B��AAu�A�р@�0A��?E_ BKjrB-5�A1��@_��@��A�G?��Z@�e�@�t@-r?ə�>���B��A"�BXJ�@�݀AX �@���@���    @�q�@k: @Ԅ@��?��?Mw�=��     @A�    >�h@^`?{��        >�g�A�z�@���@�@��>B�F?��@�@e?��@A��@v`?!��@��>��A���                                                                                                                                                                                                                L       parents[$l#L       q���                                                           	   	   
   
                                                                                                                                   !   !   "   "   #   #   $   $   %   %   '   '   )   )   *   *   +   +   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <L       right_children[$l#L       q               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <����   >   @   B   D   F   H   J����   L����   N   P   R��������   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       q�Kpj?A��.$����$>�p7��Q��4�?���I�'?���?n��?7��>� |>���>� b�W����>G�nwI?�Y�@��=��!?�wP���<?.˿.�?*%j�� ��^�?��f�d��G䓾�[&?v��xV�8��>�8��W���[Aj��~�V6� RҿN��?�b�?U�v>�>�3��P����]��?�s�s�<Ւ����>0���4�D��[��6�����˿ hL���>^½;כA>�;	>^l �cK�>���=� ���>3芾����	��*�P>�r>��f>�~�=�(�/�
<0�Žѳu>X�8�?�<Yn��=���X����^�>�$˾Dʧ;'�u>j�����)=gT��0s>/y[�5�=Wt#�<��=#��=�<^�׾C�U����>�z�;X���sǾBح<bo�>/��0������L1�>&5h�$_�L       split_indices[$l#L       q                                                                                                                                                                                                                                                                                                                                                                                                                     L       
split_type[$U#L       q                                                                                                                 L       sum_hessian[$d#L       qER�DDs��E�DT��B��JD�4�D��vDI:�B;ёB\y(B���C�#DE��C��Dl4D=
/BCBV�A-�%B�~A��TA��IB8=�C���B�)*C���C���CE�C	�ZC��D'@�B7[�D1�sAy��B��@��A�qaA�x@	*�A��?�D6A2VA,�A���?�h[?�f�B0b�C�YB��A��Bh��C�N`Cv�B�݀CY%	Bg�LB���B�AA+��CcuCi�B	gA7��D!��B�@�AW��A+[�A�m^@L�?ە�A]�A��\@6_�@��A��A|6A�?��@�_<@�i�A���@��B'&@&�Ac�CzqA�}�A��d@�M�?�X�A�aBF�Cn�Cf-�@$�Cf1A��BJ�,@#dCV��A���A��B`�BQ��B��}?��@�#@���@��2C��A�e>B�:�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       113L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       m�䢁?C��k�<EӶ?>a~�]M>���1>��Y>��M?JO!����Ka?%rоf��>��;��>d6�?D�|�j��?Y?1��?O�F�����>��*�$�??�⾘<�4ܿ_{���?�߿�ɽ��?'Cc�&ܞ?K���款m'>�ME>n�?%g�>�*4?L6Z�ƕ��g�>H�@��K?|߾P��>�M��	T+>�a�?QwV��J>��羧
�>�L�>?Ot���E?1�T>��� ��S�>��+��Z}>�b�?Z���y?;��=�9?Pyȿ+>c���|�>��@?!7��U?4^!>���?�1����_\�
;�>��V��?\!��͗�����lÿV�?AX���_3?3xþ_9?X��ʼ��>�?[�ޥ?Z��>�$���Q?U�K���>�'T>�f��L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       m                                                       L       idiL       left_children[$l#L       m               	                                    !   #   %   '   )   +����   -   /   1   3   5   7   9����   ;   =   ?   A   C   E   G����   I   K   M   O   Q����   S   U   W   Y   [   ]   _   a   c   e����   g   i   k��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       mD3�C�hB�	4B�)A�� A�=�BT�AAi�AI�A�p?}� @�r@A�cA>90A|B?���?+�Ael@By�@/	�?8 @M�@    ?� @�k�A$.@H��@8�P@�TA�q    >�*>\z@>��?A��?�%`@���?��    @�M@m�?Տ�?�`@�hL    >5� @҅�@u�?�� @�\�@P�.?�Վ?�� @��?{D@    ?��^@l��A<��                                                                                                                                                                                                        L       parents[$l#L       m���                                                           	   	   
   
                                                                                                                             !   !   "   "   #   #   $   $   %   %   '   '   (   (   )   )   *   *   +   +   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   8   8   9   9   :   :L       right_children[$l#L       m               
                                     "   $   &   (   *   ,����   .   0   2   4   6   8   :����   <   >   @   B   D   F   H����   J   L   N   P   R����   T   V   X   Z   \   ^   `   b   d   f����   h   j   l��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       m�d��.$�?��6y޿K��?���>�C�W��>�Uϼ��$��<X>�M|=�W5?�0?+0�,�>c5�Sԭ��y�����o��>~|>x��?od���@�X��	P?(,t?�@�P�վ9?a�Jm��E:���v�q�g>ŵ^?��Z�K�<��{5�%����ҿpR��;f��F�>u�JA���>^����4��?���?�⸽�b�>��v?y/ξ2��?�xh?��R?���=e�����>U*e=4��@뽫�9=�����>
;>��.���|>a<-qx>z+��- {=�����^>�Z>AvN�3>Xp�=�e0>5����s�??<�%�=�Hξ0}> (��]��\�4���.g�>h���r>>W]��"rE>�B�<&|���>5���/->�:V> |M�.�b>�.-��k=���>py�:L       split_indices[$l#L       m                                                                                                                                                                                                                                                                                                                                                                                                          L       
split_type[$U#L       m                                                                                                             L       sum_hessian[$d#L       mE;}D�|�D�}�C�5�Do�fD��C�݄C�bC)�iB��DZ�D��JCH.�B�ntC&��A8��C<$B�&gB�$kB0��B+�xC�KD4��D��B�$ Bl��C�IB�Y�A8�8B��BB�Y@FD�A�C�5@T;�B�B3��B��?�hWA�"Al�(@j�hB�QB>_pB̈�D���B��&A�$�Bn��B��A���@_�C	�2A��B�V"@��@bɁB$�~Bo ?�s?�w8@ފ0?�lzC�2@� m?�g�?��A��A��B!�\@���@�LB���A���AH��@	�-AJ(\?��B?ֶ�B ��@�e�B&�@�M�Dwd?B�cA�MB��A@T�@���A��BK�T@��BB	DA�G�@��@	��?��RB���B8�AJyB@V�NB�FA
&�@M�?��B
�_@�8�B@��A8�|L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       109L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       U;�����>���F��2��Π>�����8
�����>�*a?7|#�T	?(�v�1h>ݔ0��~�k򾱈�>�� �HX2>�Y>M@�?<�G�����⓾��>�.����?������<���
V?�\�r#=��=�x5?L������>��>�X?=>H��(�>��?�?H�4��`�>!ߵ� ;>�q�	&P?D�D��lH?JQ@��"�D���3����?Va9�ƿk��K;6�S?F�>�A���K3>��?aW?��W?1�>b|x?TD0��E�>�,$?�#?N�J���>��?	�F�ڔ�>���?55S?K�?P��L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       U                                           L       idiL       left_children[$l#L       U         ����      	                        ����            !   #   %   '   )   +   -����   /   1   3����   5   7����   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S��������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       UD51�@�� C#p    AEY
A��B�f�@e��@���@mA�@��B��m@�z�=�^     @o�@C�x>�'�@��@Wl@�QA�Aփ`@&�L@�M     >�8?�E@t�    @7��>��     ?��4?BF>.ɠ@���?�f}<�� A	Ǆ@��LA�[X?���?�f@)�@���@$�                                                                                                                                                         L       parents[$l#L       U���                                                     	   	   
   
                                                                                                               !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .L       right_children[$l#L       U         ����      
                        ����             "   $   &   (   *   ,   .����   0   2   4����   6   8����   :   <   >   @   B   D   F   H   J   L   N   P   R   T��������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       U���1<��P��n�>7!�
A�?N��?C?���?2��>�ΐ���/�%���z���>J��>���>�q@0}�?x���"*�>?��?oh?Cd��H�J�?��>��P��xP>�Ӭ��i�'�@.μ���۾��� g?Υ����(?�A^?|�l?ﬄ@��ĽP?��J?V��JA>�p7>����m^=B?���p>	'��$�`>k��@�>r��>�\�k��8n>��>���8���<���sਾ6m�>m�%=��c��'
=�
�>�4Y�e�>Uw�=��H>~�:���*> ��>-��>w獾7K:=�>%=��&=��>Ys1>?'�>zK*L       split_indices[$l#L       U                                                                                                                                                                                                                                                                                                               L       
split_type[$U#L       U                                                                                     L       sum_hessian[$d#L       UE?{�D���D�+�D���C!Y�C:�D��)B� �Bo%C
|B>&bDR��DF��B�*�?��eB3��Am�B�h@A�?lA���A�{�CR �DY�A�JD?�>B�k@�E�A��!A���@#AH�@B�4?��A�'/@�`�Al�0A �A�f@�WC�SBhݍC��CM.�@��NA��CB[D��@A�A?��|A���?�i8AuLJ@��C?�G�A2TMBߣg@"Y�AG@A@K�?�D�AFA�@}4@��k@~3�A*P�@��
?�%y@�ͺC.@�ēB,n>Aq�<B�
C��pBq	�C�=@�}&?���A��@��Bbg7B�QB�KgC��tL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       85L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       y;���?~��z�?*�.�����Z�����?5�l��<�>g�8��?T>1f��J���7~���??�=��ؾ�l�>Ď>�<$�Z�c���/�_*>�b �
�>�t߿�e��g��w��*��ܨ?CL=˹?d4�"��˿	�j? �0�?��>	���ޢ=��K��8Q>��r����h�?�������x�<�l�?(�U�ڴ��o�G���>C�B���Z�2�=&���К���<���C>�	N?G�>�Կ�?40���>���Z=��A�T,��	����4!?5��?(h���4+��� >�x�=btI�4����L>�ǿ^��ʟ����8?9�꽬C��K?�{�Ԗ�=������b<�_�����?M����)=�.K��t�=��md>.�¿E��Cz?&:Ծ/�i����A��+?�\��w�<�Jɿ_|>�4q�A���
����L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       y                                                             L       idiL       left_children[$l#L       y               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K����   M   O   Q   S   U   W   Y����   [   ]   _   a   c   e   g   i   k   m   o   q   s����   u   w����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       yCڰ]Bn�C��A�� A?�YB�`�A1��A��@���@���?
A�B���A�c�A�@W� @ƪ�@�5k?�Ւ@c��?�"T?��8?�S�>���B;�@)^@��@���A��@c@=�` AO5�@8	 @Z3�@��@��V?�e1>���?S1�    ?�z�?���>��?Ɵ�?I��?��>�נ    A�PA)�"@@��>�р@o�?d��@J$�?NۀAF��@�?n�@F=?I�    Aa]?�X@                                                                                                                                                                                                                                        L       parents[$l#L       y���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   =   =   >   >L       right_children[$l#L       y               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L����   N   P   R   T   V   X   Z����   \   ^   `   b   d   f   h   j   l   n   p   r   t����   v   x����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       y�Kpj?K�^�.$����$>�p7?^�4�?���C!�?��r?n��?=�;�o��>����d�?�����>G�W��?�Y�=��E=���?U�v��P>8� ���;Đx>�˘��^�?��f� hL��ÿW��>�q@P0�8��>�.��l+��[�:�@��?�=?�b�?!^��a�:���<��E�?�?��\�]��>��z?��ĿC!����T#t�D��?.WK;=>d���U�FY�=�2?'~�=�>8�>o��=�<��.��>X:��=�6н��<�k�-1Ϻ��t�4�<��q�>Y�>J��>���J�=���<��_���o�>px�3>\��&� �>^�M�η��)L�>3�a���<�Jҽ��S�4��;ǥL����?yQ>v�;��|2<�Z�=R%�c�3��E=Q��4����`>Gy̽S*���=����4>5�վ �1;��X�,/=ΥU�'��9��;�L       split_indices[$l#L       y                                                                                                                                                                                                                                                                                                                                                                                                                                                L       
split_type[$U#L       y                                                                                                                         L       sum_hessian[$d#L       yE@ �Di(E�#DN'�B�2�D�F�D�3gDC-�B/�BLHCBbKD@]C���C}��DF��D7#�B@�jA�EAe�B	�7A�^A�[B��D�XC\B 2C���C�4B��Cޘ�C�P0D3vAk}�A{^�B��A�Y�AP�rA8�d@1uA�F_A=�A�%@��As��@y;=B�?�� C׸�C?k|A�7�B��*A���@�y�Br"�CehSB_�~B�u)B՟�A#�_A1p�C�lB6�JC�r�B.~.D(�A&d�@�1�Ag)Z?��5A1i�A��tA>�@�,�?���A<��?��"A#�`A���?��{@��w@���?�h�A�@fo^@ex�A�@�R�?ɤ�@h�?��VBSC��IA�:�B���B�%aAS�=A�R[A�~B�J�A��2@?@@���B�A��C?�_Cdc�A��A��BLB*�B��.A��@���@�
�@?��A��A�JA���C	�,C'*�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       121L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       m�*�>��t��m�<�;�?"�οq>�;����>���=�a5?+����)�i�>�:��<�>�#ǿ=�?'<y>4����v?�W?Y�?1%Z�.d��:�>��I��?.�,u6�wj	�l6��o?�ֿRڽ���>�R�?<5��?���8��?+��>	�?![R?y1=��O?g5?3k=k�j�s�-��@>��d�(�2�GH��i�>��`?Mj7���x>E/�	�[>�dc>5��ǂv?Z�>"�8��jU�>�@Ͼڟ�>d��?8]f�s��?
�?vk�ƫ��#>�B����>��&>���?7z�>��M?0����n?(C>��\?1w2��j���>M�:�!� ��4b��RW?���?#N��֕Z?JY��o����?ǥ�����ȃ=F�&>��[�������?<�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       m                                                       L       idi	L       left_children[$l#L       m               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;����   =   ?   A   C   E����   G   I   K����   M   O   Q   S   U��������   W   Y   [   ]   _   a   c   e����   g   i����   k������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       mC��=B���B�%>Bj�Ap�`A`B�|A8\Ap@�y�@X @�� A��A��?5`?���?��?/Y�A	�@d|?=�@V&�=�0 ?� @�6h@�#�@7�`@K��@�$d@vy    >ȝ�>BP>�: ?!Z?�Q$    @T_?�]�?��H    ?r��>r�?�H�@�ڈ?�b0        >� A��>Lr�@�2�@#�r@s�?��@@��b    @-Q@�+z    ?`)�                                                                                                                                                                                                L       parents[$l#L       m���                                                           	   	   
   
                                                                                                                                   !   !   "   "   #   #   %   %   &   &   '   '   )   )   *   *   +   +   ,   ,   -   -   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   9   9   :   :   <   <L       right_children[$l#L       m               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <����   >   @   B   D   F����   H   J   L����   N   P   R   T   V��������   X   Z   \   ^   `   b   d   f����   h   j����   l������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       m�d��.$�?��6y޿a�Z?���?+0�W���Sԭ>��6�ڽ��D=�W5?�V>�C�,�>c5��n>��?��;�l�?(��a��PT>[�~�X����r?�-Q>N�}?�@�-N��Jm��E:���v�q�g>ŵ^>a�X?��Z��y�����>N?��Y��m���>�8�=�Kj>WMQ<�P?�`��,,�?n0��?��˾� g?T^?9��>vv?�w�>�Y��%�?�xh=Z\���i[><� =)\
�5w ����=����,�=�&�>]<ὒS>>�g>>'���f��]U=?�P��>)=�o>\->�>S6F���>>�=�'�>T�p�5���;=w�'��0���Xv��#�>=>Q���7>C�� �>+�Ҿ0B콬wj>1U������j<n��> �Ѿǽ��>b��L       split_indices[$l#L       m                                                                                                                                                                                                                                                                                                                                                                                                        L       
split_type[$U#L       m                                                                                                             L       sum_hessian[$d#L       mE"R�D���D��CC��DS�DD��C��(Cr�CP�BTDF��Dm�C2`�CE�/B}ԈA4h�B�XB�B��_B3�A��B�D,U�DW��C�_Bc?�B�!�B�IB�JA$.BT�@A!�A @B��@J#�A���BL�\B)vXB�eBL@x�@��0A^0�B�KA�CB���D6?�#nDW1OB���B���B�(A�u�Am�_B�d>B���BI��B*�B0iI@�"�@^s?�j?�ٖ@���?��2B� e@�ir?�_A?��ZAjx�A��.B�@�&"B�%?�h
A�Q-A��?Ì[@3�2@���AG~A�9<Bf��@���A(`A��%B@>�DM(5B ��B�A�B���@ T@q��B	f�A�*@\*A��@��IB��AA�_�B`��A��A��AR��B�A:��@Zq?�1JL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       109L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       ];@�¿��>�}C������>b?�&��=4yl���뢾fa�>��>��?+������������]�>�k���E=ǉ���>�hS����?
��>ݦ?/�����?�q��������>-~�:2w1��p����>嫌���A���m�>���gx>�j>��?" 8�{p�?g>�R�?&��>�V6���|>�r?1N�=�K��!w��>��q�5�&�j���a�?O������e@>�ǿ���p�>ѫ��J�>�wR�����\?KG��\jֽ^+�>�Z�?)?�>�����O{?,�Y<��Z?If��q>�U~�=E�?*�)>8�?l��#��?��?��?4�oL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       ]                                               L       idi
L       left_children[$l#L       ]               	         ����                  ����         !   #   %   '   )   +   -   /   1   3   5������������   7��������   9   ;����   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W����   Y   [��������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       ]C���@��@B�?> @��BO��AC� <)      =�U @=�A³UB��Aex�?ך     @7O=v >�WP@I��?�a�@8��ARA�cAq`@ώ�@f`�?�B�?�}�            >d��        @n�?%O�    @��?�k @n>�@A��@{f�<� ?�
dA��?�6`@�x?�bl@Z�?��?��,    ?��d>��                                                                                                                                                         L       parents[$l#L       ]���                                                     	   	   
   
                                                                                                                 #   #   $   $   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   5   5   6   6L       right_children[$l#L       ]               
         ����                  ����          "   $   &   (   *   ,   .   0   2   4   6������������   8��������   :   <����   >   @   B   D   F   H   J   L   N   P   R   T   V   X����   Z   \��������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       ]��D�<��P>��о���
A�<�h�=��@-F�<X�����?2��>�L��[�D�/�*�G[�4�о��4?���>��P�ֲ*>�q?iA|�q!?M5�?�	?�,p?��J�IF��c��+>3}��4�׿]�����=P1�>���>�Ӭ���'��+�K@�e�L��=N�?��x�H- ?�Y�@��I������j�.?R����&/>޵G>mf#<�����()��g�=К�ZN������(>9,��6۽�FM=6&��(�Ǻ�=����rmb=�0�+����Ӣ>s�@��M~>
6�>KX=�Ʊ��>O�<�j>qT��ջ> �c W>L�e='�>4�O�D_[>-h�>2<�>YL       split_indices[$l#L       ]                                                                                                                                                                                                                                                                                                                                             L       
split_type[$U#L       ]                                                                                             L       sum_hessian[$d#L       ]E)>�Dz�RD�@DY�CZoDn�KD;Z5DX�?�_�B��BY�VC��vD%�CA��D
ݼDT�TA{��B�X@[�dB$B�AU�OC!�|C�oB���DQ�BR�iCF�B	�DA�Ahޡ?�oB���@-�'@�?�n�A�<�At�i?�YA8��C�PA�Y`B= MB� �BϐA$޵C�sC�B(\bA)DB5}fB��dBH?΀�@�>D C�?�Þ?؞�A=/nA_J2A��@�??���A"��B�3�A̜gAt�A]��B&��@���AV��B�+�Bqw@k��@���@��CcC��CF"A\��BG@�@�@:lU@�RA�uB��?�yB���A	�A�K@a3e@�|�BxF`C�~�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       93L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       k;��D>�p�Z�?(]�;���>��)�?_���Z>`Z��JK=��Ͼ�������2A?+��>�|=Oł�>� ���C��}�=S>��\���e���!ž�7�	��q���u>���?3D�?� ���־05�>��?)��>^,c>m��Ҿ��?�۞���a?�b>�~�#
w�SQ�	%�̶��A���	�c#���=}F��Ƃ��
���>Y��>I�L>ǁ�%?4-�=��?'�b����x��=����P���3q?��?;��>��"��Դ>�;�?"���C9�*�>�f2�;�����?U�4�>.���C�>E4O��6˾�������+Z>�E�I��� ⨾�=�?�N���6�n�>�w��������=4�?UG���Mؿ8��WkL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       k                                                      L       idiL       left_children[$l#L       k               	                                    !   #����   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q������������   S   U   W   Y   [   ]   _����   a   c   e��������   g����   i����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       kC��tB>>�B��LA��8A_�)BO�]A$��A'�`@N\.@��u?r��Bf.�?��@A!��@D @���A$�@ia�    @ ��@ܗ?���?��B��AN,�@��>�� AR�?!
`@���?&� @G�V?�� @�P?��t?��?	�(>�@ ]?�ۖ>4�@?^{l            A`WPA��@��K?=�@��}>2-`@
��    ?j��A���?�Jr        @��"    ?�                                                                                                                                                                                         L       parents[$l#L       k���                                                           	   	   
   
                                                                                                                                   !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   -   -   .   .   /   /   0   0   1   1   2   2   3   3   5   5   6   6   7   7   :   :   <   <L       right_children[$l#L       k               
                                     "   $����   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R������������   T   V   X   Z   \   ^   `����   b   d   f��������   h����   j����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       k�E�/?��.$����$>�7l?=�;>���?v�?�Y�?��"��>��о��>�������W��=9F�C!��0m��o�쾓'�0S<>�5��>*��d�>��z�D���;H��v�BH�?|� @AH@�@�V>�,���[�O=W��g,@S�P���Sw�5��a�>.�>�8�?�j>��e?|�G�]������>ﳂ�4v����~>�Y����2�پ/W?u<="X��QB=�g��1�`>X7<��>Hi齇������*y�=����`߼�
�>.�$>a-n=��)���=��>C!���#�L�彊�aC��(��>Ϛ�(?V=Q�B���=l�,��A���,�4�=�(4=���r
;A��X(>6?+��a��$=�)����3<Xm>�]j�1��g�L       split_indices[$l#L       k                                                                                                                                                                                                                                                                                                                                                                                               L       
split_type[$U#L       k                                                                                                           L       sum_hessian[$d#L       kE*Q�D[dD���D6C$C��Dt�DY��D+�B2�]B��B~k*DH��C,��C���DX�Dq~B�:{B��AwB�A]��Bk�Y@�n�D�RCW��B��C�C=�B�_�B"[�D3"B8��D�cBz%�B O*A�_�A3��A��|B[�s@��A4YBYAͼ @#D@��C�e�Cf�B���C dMA��"Al�B��B��B�8�B���A��RB�s�A˳�Ar)?��bD�]B-ʫ@.q(D�@L��Bb��@�~�B`p@�u�A$��AV4i?�ՄA�DAD�4@t7AM�HB(@�@8>�?Ӟ@�!U@&��A��A�WC�6 AE�C/�B�k�BT��B	C�B�KB�X�A*�nAGA�@�lAH��Br?��AЪEBL�B���B*|nA��j@�S�@�_'AX�C�G�CE.DL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       107L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       W�d�H>�bG���ѽ�@?�ݾ�$	> �&��s>cV�>y+G?��OY��.>�yl����=�X?��?� ���Z?
W?!�����B�=�s���9?s���U��?�n���>ʫ���"=Fhh?�X��sB>㒭>�{�? �p���'Bn���Ŀ1�>yh���I� �?=�x^>¤�?8)�K P>���� U2>�1
�Co�>�*���y�)߾}v�?F->��2?'1m����?{ъ?Sv��_>������ݾ���>�u���>wǪ<]L�J6=V��?^�	M��r���z�)?\<P���l?��=�gE��xn>�lS?�Y���w�}�+?+�1L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       W                                            L       idiL       left_children[$l#L       W               	      ����                        ����      !   #����   %   '   )   +   -   /   1����   3   5   7   9   ;   =   ?��������   A   C   E   G   I   K   M   O����   Q   S����   U������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       WC�R�BY� B���A�rBA�:�AlD�A�@�    @�a3A��V?N� ?��A�[A\�??��@��    ?�� AO�@"[�    ?rB @b@�9@<O�@0*�@���?�    @��>���?cY>D��@�{�?�c�@UD        ?���?҄>�#@@���?�|�?���@F]q@�*�    @5{-@���    ?�                                                                                                                                                L       parents[$l#L       W���                                                     	   	   
   
                                                                                                                       !   !   "   "   #   #   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   /   /   0   0   2   2L       right_children[$l#L       W               
      ����                        ����       "   $����   &   (   *   ,   .   0   2����   4   6   8   :   <   >   @��������   B   D   F   H   J   L   N   P����   R   T����   V������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       W�d��A��?��� g�.$�=��E?+0�+|$>�8��Sԭ��<X>�M|<�h�?�V>�C�6[�>2����P>��;>~|>A�@���rW>f�
@�u?�-Q?��~?�@�#�ÿo�>��[3>Y~R���?���?q�u�F�>A"�.a�����>�J �+�K�քh@E�]�������>\�@`]>�-:���?�xh�j�]=�̚��+�,���>��>��>H����3�>�S>�[���?> �-�����e>����=�� ;��Ⱦ#�A<��.>.q�$Ú���� �1F>�$0��?�>=�<�{���=�1>0K8��r���c�>NcL       split_indices[$l#L       W                                                                                                                                                                                                                                                                                                                         L       
split_type[$U#L       W                                                                                       L       sum_hessian[$d#L       WE	�Dr��D�:�C�=DK�7Dy�Ck6B���B�0�C8R�D��D26qC��LC7ؕBMu�B�
A�� B�тB�ӚB�Q�DPVD'=�B/�\BđAC;}�BӋ�B�%]A��B)�NBg��@�)L@���B���B�sB��B��B�}D%�t@�;�A?v�A�U>B���AÙ�C2zA��Bt{B3BPmXAϺ�@��c@U#wAi@B-l�?�l@��1@A�?�24B
R�B5�BxЎ?���B�@<<~A�@�Q@��?�J�@qY�A |?�{�A��B<u�AտRA���@��C({A��@MB@��BNPA�|UB5�@�rA�� @�Ҕ?�!�?�%>L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       87L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       Y;T4���>��	�������=�i?���`=&׼�����b��Զ>���>�**?����c����Y)�]�$�CR�>��ᾥ�A>9=�[>?�~�2'�>ھ�>�? �
�eh?Vi=��\�������>Z� ����?.�C�s��
y�f�>j�4���}>�>�S?n�Ƕn>��F>b��?	��>�=�]�>p8?!�k�x� �K�<�O? d�>$����=���T����=cf�e��@\���>�y��A�?99��>�o>5��?3 �?Ȑ�%Y�����B?"=8���5�>��>�Q?*[�>���?�J���>�$[���?�dL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       Y                                             L       idiL       left_children[$l#L       Y               	         ����                  ����   ����      !   #   %   '   )   +   -   /   1   3����������������   5   7   9����   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W����������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       YC��^@�� Bz��?+ @�ArBFuA�P=�h     =˳ @֐A��A���AǴ?��    @     >Y��@!8�@	*�A�A �RA���@>`@ii�@��@?�1�>�D                 ?�b�?���>�    ?��PA��@X��@��8@���@T@�g�@.c ?g��?*t�@j�@@�?u ?�t?p.�                                                                                                                                                    L       parents[$l#L       Y���                                                     	   	   
   
                                                                                                   !   !   "   "   #   #   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3L       right_children[$l#L       Y               
         ����                  ����   ����       "   $   &   (   *   ,   .   0   2   4����������������   6   8   :����   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X����������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       Y��D�<��P>��о�����?�C�>�wt@-F�<H6?���??��>�\Z�?�n�` l�RRо-vw���4�-7�?�@^?2�ʾ[>ؾ6��q!���� hv?��?��J�UB��4�"y�>"g�<�o��D�?
X��[ʽ�'�>Q˄>��P�[�:?bV�.��?Qپy�@�@i-�L�h88�A�ڿL��H�X�T��?@�&>B>�<t*�@���bG�>P=D�Ǿ�%�7(�<"�"��<!D�'G,�9��j�=�����>*��"=�R%=ZCo>V͋>=W�1�k�-���'Ń>8��<]�I���=�?I=�ǵ>Lm�=��>3����=��n��;<>(��L       split_indices[$l#L       Y                                                                                                                                                                                                                                                                                                                                  L       
split_type[$U#L       Y                                                                                         L       sum_hessian[$d#L       YEk�DJ��D�}�D-S�B��BD]�D%
D,�v?��Bz6�B[��C�4C�4C]��C�3�D)��AP�iBp(e@ ��B9��A��C\��Cn��C=�Cn�A��#C@ݼB���C�ʈA<��?�&�?�%?���B�NA/�y@>��@��BB��B�BAI�C>P_B���Bئ�B�>C#�A���A(iB�v�B�D�B�u�Ax@phC��A9!�A�=�@��/@�4�?�3�?��B�@RAMn_B�bB��A��yA�#Bz"B���B��<@�D�@z�CB���BQg�A�(�Cgn@�҉A:KoA<p@�/?@~C$@��B{�\BH$B�B'A�B0��@ �@�?�D7@��L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       89L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       i<!/>�%�lp>ܹ����`�	n��/i?w6�F��<�Rܿ@�5k��
�������?%�=O�w��_=�,v>�u����>��9�;�>����6������}�U?<�
�����9>v@�?�>�)��.�>C�z�d�>�+L��ks>��w�]��;I{��Ϧ�����&�>kJ�����4k��^���$W�
Ry��"<��ݾ�{<륝>Po� H�?ڳ;��?#�>#�~?	�־�P�>$���+$���?
�c��A��J�>�0t�۰�>�����|]>�>���ܽ��c�r
?�d�U�JAC�f">��ؿ�">��ξ��J�'>ַ >976��q^��X�d����>e{$�B�������]?? �t���'��>�m����@�?VL���B�c�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       i                                                     L       idiL       left_children[$l#L       i               	                                    !   #   %   '   )����   +   -   /   1   3   5��������   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q����   S   U   W   Y   [   ]   _����   a   c   e   g������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       iC@��B���A���B5��A�ٜA���@k��A���@���A?��@@A�͖?���@���>_h @�� A�@� @�j�A��@���    > A��B@�B?ڞ�>��@@�af        ?��@@��@�^`@� 
@[�?��*>M��@h�@ǳA	2�@d�@��?�Xx?�Z�    A<�n@&9X@,�(?��@E��> K�?ݳ�    ?~ΐA�?�^	?[�                                                                                                                                                                                                 L       parents[$l#L       i���                                                           	   	   
   
                                                                                                                       !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   -   -   .   .   /   /   0   0   1   1   2   2   3   3   5   5   6   6   7   7   8   8L       right_children[$l#L       i               
                                     "   $   &   (   *����   ,   .   0   2   4   6��������   8   :   <   >   @   B   D   F   H   J   L   N   P   R����   T   V   X   Z   \   ^   `����   b   d   f   h������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       i�6�h���.$��d�@��?=�;>� b?a�	�A(�>�7l��~6=�k%���?�0�ݑ�������Ŀm?�Y��-��>�fR>�V>�I�?�>v�,�d�>��z�/r�&:I�+�� ��5�r?Ap&@%�v�can�������K>���X��?�j?pŝ?)\�Sw�; ��4.�?�&�?�*��-��҈�]������>ﳂ�+,=�d��<{�>�q����>8�
;"t>>��=D��>%O��`�=Eͩ���_����>&��ε3�*�
>���Ѐ>��J�>?���ռル�*�@>=�}��U3�r��� )>�����=����ָ��2ܖ> �G=^BA��Tؽ�� �6�N�1]=��I�i���4���	�>�%�v�+��=؃���н�<>��M��P�#�,L       split_indices[$l#L       i                                                                                                                                                                                                                                                                                                                                                                                       L       
split_type[$U#L       i                                                                                                         L       sum_hessian[$d#L       iE�D�gD��hD[~C֟�D�bDOnDA�B�/�C� SB���C�$�C��C1D�C��}D,��B���BPT	BH�C�nB��o?�(B�5IC�z�BީlB	B⋧B�3>B�V?CU�kC�BR��D]�BИB:96@�Q�B=	�B�A�k�C*�$B�B�B*B�(�@��Bl��CscB�aB%pzB��/A���ANj�B�ZB���B8s�Be��@W�-C�A�K�Br�D�B��B�@��A)�B�?ܒ@FZfA<�B�A�@M@���?�MVAo�B�=�BP1B}IA�xA��A�VA�/5B+:?��g@��gCU�A�l�A���@�A�-9A���@���Bzd�A
��AK^�@~�A+�4A��'?���@���B��B�2A��?��7?��$A��B�J@L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       105L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       a��B(>����������>�L���+�=��S�
>�><P�>b`%?-�� ����C>�G*��Mt=_s
?PD??��j>���?�{�	w����>z�%���? ��<��>��'�/���l>��}>��n?z�=]�|?�+����>��a>oI�?S^?	�<�
@h���E�db>���ӿR���F>&��?��F#>�M��.>��=��r�������>`;־�l�>�̾� �?�־l�>��f>��\?VX��W?B!>�K��$>�CM�Ι�>�?���E����>�1��������? *��6!��ۿ1R�?%>}�{�>�?��52?"f��,��[�>-M�>�N�� M�K�I?z>8�f���L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       a                                                 L       idiL       left_children[$l#L       a               	      ����                              !   #   %����   '   )   +   -   /   1   3   5   7   9   ;����   =   ?   A   C   E   G����   I   K   M   O   Q����   S   U   W   Y   [����   ]����   _������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       aCj��B�.B]+A�gfAl��AXd�A��    @o��A5��?W� @qU�A6$KAȅ?M� @#�=eB ?_� A��@     @@@�v�@�i2@`z$?�N�@���?�H�=�� @p�[@�2?�˪    ?I�>�� @=t�?��@'�v?�V     ?+b @�F�>�\�@)E�> �`    @hK@��?iI�@^52@��|    >��$    >��b                                                                                                                                                                        L       parents[$l#L       a���                                                     	   	   
   
                                                                                                                           !   !   "   "   #   #   $   $   %   %   &   &   (   (   )   )   *   *   +   +   ,   ,   .   .   /   /   0   0   1   1   2   2   4   4   6   6L       right_children[$l#L       a               
      ����                               "   $   &����   (   *   ,   .   0   2   4   6   8   :   <����   >   @   B   D   F   H����   J   L   N   P   R����   T   V   X   Z   \����   ^����   `������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       a�d��?��?��� g�.$�?��z?+0�%�>�8��Sԭ>~|���D=�W5>���>�C�`S�% '��P>Fz:��~>7a�T�>[�~?q�"��b�?(,t>��?�@@�9<lgA�����k� >.�9>Y~R>0+?�Y�?gyg�ER�㳱>%�?�`��,,�?�ֽ%����'�!/Ҿ��>��v@<F?�w�?���O?�xh�$R�?hr���Tw=��N���>��4>'h����>�
>�k>;�н���>h�(>:����&=��]����=<^ >5
��(�S��BL=(�n�R¾,�x��ne>�żZ��8�ԾT��>FJ����=���"?�>4)H�N$���e=O�%=�+����tE�>=��=]��X�L       split_indices[$l#L       a                                                                                                                                                                                                                                                                                                                                                           L       
split_type[$U#L       a                                                                                                 L       sum_hessian[$d#L       aD���DK�gD�C
��D)CDOM�CS1�BS�B�a^C%E\C���D/v7B��'C)�KB$�B{�A�{�B���B���C9�C��D��B��2B9�IB��B��yB�@��bBUB)�zA�z�@�
_A���@��B��Ba��B7�A�oB�ъ?�K�DQKBf��B��?B(a�@��BO� A� 	Ab��B���B/mB*��@�߻@H;OA��@��~A�?,A�O�@ZOA�7�?��@�=@:�?�B��B'�BZ�
?�CA��@K��A��@��gA$BϮ�D�$B"}A��zA��SBM��A��3A�T�AD�_?��L@IN�@�nCA�dxA2Tw@@�B�]�?�(@A�m�A���B�@Ҫ|?��?���?�˓@aq2L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       97L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       Y;L�#��&>xDп
�;�Z=��>�l��Rp=&�s�����eO�v�><-�>��|?F� g��2A�9*+���U��>Ot־�S�=�m;��H>q��=o��>� �>�g�?2}�v>����j=�F쾧`�>�rL>��X���׿c��+���x0�>yJ���s>��]>z>�����?�>��?�f>��=�>�U?6����r>�R?Gc�<Ѿ�~l>�k��6��������>mu�̃?>r&>�uI��JC�e�g�L?PR�0�����>L�Z>�%�?�ξ�M�=1Ɉ=�d�?-͠���>��>���?,u>��?�����>Fi�6?�)L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       Y                                             L       idiL       left_children[$l#L       Y               	         ����                  ����      ����   !   #   %   '   )   +   -   /   1   3����������������   5   7   9����   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W����������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       YCy@�@��@B1a>�� @�ҘAƠ,@��>�     >1� ?��AI�A���@�T�?Ð�    ?�E>-��    @%�?���@<�@O�)@�aA&�8@�ī@3�?���>ɲ                 ?;�?�К?��X    =� @�?�A�@&�?�0?�7�A2�@O1 @t�?V}@@�h?Ԯ�?U��?��?�8�                                                                                                                                                    L       parents[$l#L       Y���                                                     	   	   
   
                                                                                                   !   !   "   "   #   #   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3L       right_children[$l#L       Y               
         ����                  ����       ����   "   $   &   (   *   ,   .   0   2   4����������������   6   8   :����   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X����������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       Y��D�<��P>��о����Ҿ,�>�-z@-F�<HM���jt���P?E�v�[�D�%;��RRо(&���4�V��'�x?7�޾��>�ΐ�M�?M5�?y}@�?��J�UB��+���Z�>j��8�<͈O@4]�������'�� e?2ڼ�a<?��-?��a=N�?��x�@��$r��<�v>�q��L��H�X�T��?�R>3=��F�=�w�>oD�; �.��1O>@��+ۓ��?��
�=4�Z��jL=�J	=��%��Y�F
���><�ɼSY��P�=uݠ=ȓ�>8̑��*<UX==o�>P�Z��%�=��=�^(><��=�3 >"��=�*?�Zz�>4��L       split_indices[$l#L       Y                                                                                                                                                                                                                                                                                                                               L       
split_type[$U#L       Y                                                                                         L       sum_hessian[$d#L       YD��D"�MD�{�D	,B�9DL$D��D��?��BGNnBO#�C.�D fCQ �C�'yDMA-��@'�NB<��BٹA]'�B�B���Bp�,DY�B��!C	��B��C��A�?�Vt?��G?��TA���@�#pA:��@
�B�_A��0A��mB<Y�BE�A,�eC��yCJPB`#�As��B[TB���Bba|A'�A&�C�k�A�<?�u�@>�@���?�-A"�+B�-�@��A��SAJ9�A^��@���B'uk@�"}B1y@���@�H�@�O�B0~�C�{�C&B�T/Ay8tB!�g@�,A3_�@���BEC�A�ҜB}h�A��|B�>@N[@̨V@�s@���L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       89L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       e<Cg>q�3��}9>�Uh�DG���M���t>��˾�c�<���N���醿��������?x> ��^�>�T=�UP���b>&|�'�=�~��k�<�y��S��GJJ�	� =�����N=��#?��>w�7��<��i���_>���*�>sH���/>�Z��lؾT�t���>xAw�K������bq>���S���Ye>����=�>��m������G���>�rU�uO�?8�>�)>�-X���.����I��k�>�p\?-'��F�?j���q����>�q���7�����(��?���)��>Ӯ����H��Z�>�e�:��۾��$>8dL���=B�i�Ͼ�M�>��>.����)?�f���,>�ݟ�<�Q����L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       e                                                   L       idiL       left_children[$l#L       e               	                                    !   #   %   '   )����   +   -   /   1   3   5����   7   9   ;   =   ?   A   C����   E   G   I   K   M   O   Q����   S   U   W   Y   [��������   ]��������   _   a   c����������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       eC|�B>4AǹA�qHAS�A�[�@_B�At.�@���A�i?D<`A�f�@/H ?�@��A*�0A !�>��?�A�@ļ    >���AM��@�P^?��>T$�?��"    @Sx?��@��o@*� @�P�?#�?���    ?�?�?펄@؅ @O7�>��?`�8?� ~    @��@+�c@%��>�* ?���        >Ы�        @w��?
�\@$/(                                                                                                                                                                            L       parents[$l#L       e���                                                           	   	   
   
                                                                                                                             !   !   "   "   #   #   %   %   &   &   '   '   (   (   )   )   *   *   +   +   -   -   .   .   /   /   0   0   1   1   4   4   7   7   8   8   9   9L       right_children[$l#L       e               
                                     "   $   &   (   *����   ,   .   0   2   4   6����   8   :   <   >   @   B   D����   F   H   J   L   N   P   R����   T   V   X   Z   \��������   ^��������   `   b   d����������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       e�5n���.$�>�R�@	�?��ʿd�>�ٴ;=>d��A��q�>/�e�� hL�쿃�?!D��Y߿k�?�c����=G�>�I�>�}>v�,@hr@S��FY�%��?'~�>�Vn>&An>� �@�?R���^�>�,I?>`^�>��b�V�r�#v���-�?b��; ��,48���b��V2�t�ܿ@�C�1���5"�?n�=ʺ����/����̦>�I��(�9=��/�>3�=�ܘ=�����Q�ľ$%�@�=�S�>O����*>����w���6=��{��ܽ���J�y>+�9����,o�=�(��_��r=��9�n���,=]E)���i<i�K�,�ƽ�]}>d=Q�Ľ�We>V����=/;��=&�bJb�p�L       split_indices[$l#L       e                                                                                                                                                                                                                                                                                                                                                                         L       
split_type[$U#L       e                                                                                                     L       sum_hessian[$d#L       eE��D���Dg	�D=�kC��rC�ƆC�L�D/��Bc{C��;BR)�CȤB��CY��C\��D}�C ��B�A��C�{�B@b?��WBM;�C�l0B��HA3�B���@�ICS�B�OC8��B�G!C�i>BӍ�A��	@�a?Bt�@�KEA!C,�8B�y@R�B3A�@���B7�sCG�B�{>B,�&Bu6k@��@A�B��"@{.?�Q�@���A�R�A�B��QB� �B1G�A���C�{B^�B���A}O�A��AY&O@o�"?��@���?���@A@��A��8C��B�)B��?�=�@	�A��A��*?��k@~�AğC.��BҦBg#�A�ZYA���?���Bq)K?���@�&_?��x@5�bA���@�7?�۲A	�UBQf)Bv6zL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       101L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       e��!>>��\��H����>쿈���f=�nx��=��>s��?QL���+�F� >`�{��\k���8>�S���e�>�h>�Q?��(f�9�I=h�S�䊯>�SA<�{t�I����Ⱦ�[�>G�>>���>:�οdi>[�*?�>vR�?�q>ݿ5?4=�IؼJ u?
X��!8>ɪ����W>�����>��|?����p>�/>b`[��GԿ	��=צ�?7�� Fm>�1����>�>��T� �?�<���?��?���k6�î>�b�=[E�?(�>�S��V�z���?���A.?.RB�](>�F,���?&3>���K��?2�}�6	P?MD���@��e=G�x>�z?�g>������Y=�*D?ʚ��!0=�g��/TL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       e                                                   L       idiL       left_children[$l#L       e               	      ����                              !   #   %   '   )   +   -   /   1   3����   5   7   9   ;   =   ?����   A   C   E   G   I����   K   M   O   Q   S   U   W   Y   [   ]   _   a����   c����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       eC$�(A��BW��@��<@�`A@Y�A��    ?�)q@���?���@-/�A1I<A�b>\��?�b�?'�@+�X@(�x?���=�� @��@~u�@��@�?�İ@��O    ?mQ8@�<?��?ũ�<�m@?�D�    @��T?��@��j>X|@?g@    >�� @(8?�?��?��@� ?���?���@f>Yq�@���@��`    >� x                                                                                                                                                                                        L       parents[$l#L       e���                                                     	   	   
   
                                                                                                                                   !   !   #   #   $   $   %   %   &   &   '   '   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   6   6L       right_children[$l#L       e               
      ����                               "   $   &   (   *   ,   .   0   2   4����   6   8   :   <   >   @����   B   D   F   H   J����   L   N   P   R   T   V   X   Z   \   ^   `   b����   d����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       e�P7�W��>��.�� g� �*>�dL??�ȾM_;�lླ���U?�#S>�3_>fw�?�V�^�W���T�>w{`�F̾㳱?O�⾭�оˈ��n?(,t?� �#��?��J��[&�`qS�|a��l+>Y~R�"x~>΀?��f>7H0�x'����j>.>��4�>m<��Qؿr���Վ>*X罿�6>�̏�Hq�?y/�?���?�~�=��j>�q�%��=d>[���=�Ռ��|�=�>�̽��>+��;��>,T�>4�ҽ���1Q8><��(>,��>�̽!�ξ&�ƾ��>#܀�'>Q/����L=�!�F=>G;�='�H�t��>VT0�Zq�>vR��ⴼ	r�<o��>�J>0.|=�� �̹8=�)>9���<�I��� L       split_indices[$l#L       e                                                                                                                                                                                                                                                                                                                                                                         L       
split_type[$U#L       e                                                                                                     L       sum_hessian[$d#L       eD��D��Dp>�B���D�D.]C�DzA���BOb�B��Cɫ�D�_C-��C]�8B*>�A�G�A�~	A�q�B�IEB��(C���C��&A֙yB��IB���B��B���A��PAS{&A�&�A:B�AT#�A �)@�"�AeRqBi5�B!]	B!*eB6w�A�3*C�tOC��A��@�mA�X^AлmBuL�@M��B��BF�nBe$�B�iJA�>@�WA3A%f�A�G@7j+AhNA^�@��4?��;@��@�a�@?�CB�A�h�B��?�IA��A���?��pB2@ A���?�:C�BB��@n<@�%X@��?�MH?��A�{\AE��A[��BZ=q@�{X?���?��)B�.�@�a�A��bA��yBJK@���B3`�B!q�AЩ�@k��?���A�`L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       101L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       W;�8���D>Vx6��꾑5�=�>�ѿ�¾���aP��k���>u�>s%>��e��`6>ѥ���2���G�F>>�!���d=Q��=U��>ȝm=ZX>3>��F?	o۾�a�=��׾�N�>��.����>��\��y꼯$=��>�q�����>d�>We>򧤾r��>N�Y>\�x?�>��>@§���?
�N���<}?4*���k?1��=�	���Hq>X�=����!]��YaE>&6�?�-��uD���>�0�=�"�>��Z=��z?��? �H�䈂�޹w=͂���y>�
�=r�s>�f7���?lS>!Z?z��4��>���>��?��L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       W                                            L       idiL       left_children[$l#L       W               	      ����                     ��������   ����      !   #   %   '   )   +   -   /   1��������   3   5����   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S����   U������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       WC3]�@��B�'><� @w�A��0A
�@    ?��>>�?�y�A3�A8�@�[d?�ۀ        >3d    ?��v?��@��~@ϟ�A5��@/�H@�v@J�(?�^@?I�         ?7�x?l�}    ?q��@/8@D�Y@��@b��@b�@�@>r@�(@$�@}+@%�y?Rc`?y9�@���    >b�                                                                                                                                                 L       parents[$l#L       W���                                                     	   	   
   
                                                                                                           "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   2   2L       right_children[$l#L       W               
      ����                     ��������   ����       "   $   &   (   *   ,   .   0   2��������   4   6����   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T����   V������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       W���<��P>���@-F����?�C�>��h�$3����4��jt���P>:�@�(�	?��J�RRо�=��k�����#*�?7�޾���?Pp?�	�	|�#�x�	T��L��\W2�<�`���<���?
X������X��u?���@:�4�@2�?Q�>m�@�@i-==)�?R4?n�X�#Kܿf��[� ��`#��-��"��b/�>X2i��8�>U�<��K�^�=�((<�ϾA����m�=Gt�>"�н���ĺ=��A<Ԑ=��<���>2��>tW�	���{<��*� ��=�ن<���>
!�-Y>/�1=A8m>,,ҾX�R=�R>��>.��L       split_indices[$l#L       W                                                                                                                                                                                                                                                                                                                               L       
split_type[$U#L       W                                                                                       L       sum_hessian[$d#L       WD�!QD�D�;BC�q*B��DD1�?D�FC��A�^BxQBC�7C���C��CT	bC�#�@�iw?��@ΓB[gB�bAO?SC�OCV�FC��C>(�B�GB�˸B�өC���?��e?���A��@ȟ3?�3�A3�Bנ�B+P C/iyBO4B2ŃBޚyBqabC�sA��Bw&Bt6$BgaLB	��A��?՗�C�XAu�A��?���@��t@D�A��B˝*@�7HB^w@��AB��UB�4�BB@�e�B'j�@5��Bl�:BP��B5X�Ap"�B��*@���A���A<��A���BܳB��A�7>@"}B]?�ASA˂)@\�A�RB�I�C2��L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       87L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       ]<j@�>X�;�pȩ>��0���r��O��v�>�ľ��="}t��$ �\���Խ��9��nl>� �S�p���=���>�}�Ap���cP���=�_S������$��'վ�Ô>�Nb���u>��=G�<<��a�
��>Da���>�>wx3��T]���n>f|�<�L��=]>� ���]���
y]���>;�ϼ�b'���F���>�`�>=���>����?��>y�>?(�о�x�?�5�BѾ��3?�ݾ�0�u�>����T>(s�ݝ�>�Wf�ͪ>����z�>��&k8>���Ç��i���
�J>����M�=�Sž����4�	�0��L��
�)?}F��sK=}4ľ�!�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       ]                                               L       idiL       left_children[$l#L       ]               	                                    !   #   %   '   )   +   -   /   1   3��������   5����   7   9   ;   =����   ?   A   C   E   G   I   K   M����������������   O   Q   S   U   W������������   Y   [������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       ]B�zjA��A�@2A��A$�LA���?a~�A%�x@rm@�f%?F#PA3	?�[�?���?��@�e @[&?��L@]�MAT~@7r�?��>� AK�}@��8?�]P        =~��    @	�@��pA��?��    ?� >��@?��D?h�@K�@��@GI~?�                 ?��A?�e?Z:�?�x            ?��?jR                                                                                                                                                 L       parents[$l#L       ]���                                                           	   	   
   
                                                                                                                       !   !   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   /   /   0   0   1   1   2   2   3   3   7   7   8   8L       right_children[$l#L       ]               
                                     "   $   &   (   *   ,   .   0   2   4��������   6����   8   :   <   >����   @   B   D   F   H   J   L   N����������������   P   R   T   V   X������������   Z   \������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       ]�5n�'��^vܾd�@	�?-M�x��?�R�A(�>�E,>�I�=��D?�ƾ�v�QB?8��=�9�m?�Y���>��p�; ��j<�����>v�,?��*�3� �������#Xu��5�� g��`g�Q�ξ&T|�X����K?*	��Wfٿ���?��r? ���U]�>z ��8��Ծ&+=���?��:>�px>�>�2>�>��<݆[?S��uv>=�ܿ>Jwa���>*=ڽh�b���q>66=��m� &�=�Ӿ2x=J#���a=����!=̞�;��>݉�G��=$5)��Ƚ�'��&��=�ֽ됈<�1S��aG�;?�%Cm���)�&�e>Ɉ���[<��v�z�L       split_indices[$l#L       ]                                                                                                                                                                                                                                                                                                                                             L       
split_type[$U#L       ]                                                                                             L       sum_hessian[$d#L       ]D�3�D|�vDG�D ��C��oD
fQCu�#D��B�ߌC�nPB)��C�HsC#^@�8Co�bD��A��B'AB+��Cb~YBļ�@��jB��C���B��B�ԤBLx.@jS�@(�C	��B�i3C�Be|Ax�WA�@�fLA���A�6AA�RB�FC<��B�Bn� ?�yZ@b�'?��BABK<�Cn�XB(<�Bk�B�I?��?���?��`@�q�B�rC�y�B�#�AU̘A��@}��A9Q�@Y�@r�A�sA�^�A�t@),�?��A01=@�/xB�WC��B\SHA9��A�-�@���BT�FA�t�A��CT�pAϧ@BMNA�@�+BM�>B�}�A�,�@i�p@�@JwB�XL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       93L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       c���	>�\O��Ȍ>
(W?�u���v=��_�,K�>�"�>��?<��*��>%И���x=������>���=��^=�ʽ>ڣ"?�>Jm��%о)�>�����;+R2>�1-�߾}�˼i�?�?�����>�Y�?V��iu>�_A>>Iþ׫�>F�>�C��v��"->����ڃ>g�O�%��?�>8n0�N_�>��8>�~q���;�NM>#vd���>@��>��-���>??�!?w�>Wܿ�+��>��8>��<��y>���fD�*3�<K쾬6�>��g�����K>�=þ��>�u\�.@e>��� d�>���	��"n��o�>�+���6��@��?k�X>T微�=?��A�)>���}R?:1Ҿ�d�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       c                                                  L       idiL       left_children[$l#L       c               	                                    !   #   %   '   )��������   +   -   /   1   3   5����   7   9��������   ;   =   ?   A   C   E   G   I����   K   M   O   Q   S   U   W   Y   [   ]   _��������   a������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       cB軯A�J�BF�A��@[ A%A)e,A*@�[�?x�<|� @	�@@��@���>�M @9�?���?�
 @7v|?�*>2/�        ?C� @+gx@b�?�5P@�,Z@�ED    ?�Tf@IW        ?��2?���=}� @-u?&�?ҋ>�B ?nqp    ;�� @k,�?3�x?�o@3jX<�o�?�*0?�@o�g@��?��        ?��                                                                                                                                                                        L       parents[$l#L       c���                                                           	   	   
   
                                                                                                               "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   8   8L       right_children[$l#L       c               
                                     "   $   &   (   *��������   ,   .   0   2   4   6����   8   :��������   <   >   @   B   D   F   H   J����   L   N   P   R   T   V   X   Z   \   ^   `��������   b������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       c�d��d�>L �����?��?���??�ȿT9x�@��>�8�=�>�8�>�3_>�<?�]�?Mo�� g��FG?��NL!�% '>+$ =r�>������?g��@�?��?�*T���?�2h�>2��� �I�*�>ŵ^������ g?��f�;f��=m��k� >5)��%��ְM>��P�)2�X�?����@;��QB?U�v@�D�6�ȕ?�����=g;�=�c�"4=e@�> h(>-\�=��s�M�l=�'�>��<��=��U��þL>	;s�O�Χ�>���C�"��=��<>y��Q=�W�Z=�q�%OV�B덾9R�=��S��g_�>�o5=~xG�ѻ�>'��h�2>��ޖc>_n����{L       split_indices[$l#L       c                                                                                                                                                                                                                                                                                                                                                                 L       
split_type[$U#L       c                                                                                                   L       sum_hessian[$d#L       cD���DP�D<58C���C�
QD��CX��B��C4��B	��Ck��C�dzB�ZJC7��B4Bq~�BW��B�_B�V�A��-A� "Cj?�S C��A��BE��BO'�B�7�B�k�A���A�BM�A��B/��A E~BX�jBx�B-=A�/`Aw�W@|
@��AC}QC�1[B�	�@��\Ad��B/$�@�BoB<
s@��>B}poB�>B���@�n�@��@`N�A��A��@�"�@�h{B�uA���Bo��@�B *GA3��A�б@b�wAT�@
yV?���?�^p?��B@G7�@³�C�&�@��B��@�a?��?��AI	�A�vAa��?�� @�Ч?�ĺB7�M@l\?�j@A�?DB=P�A�WA;N�B���@̍�?��.@�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       99L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       W;�㽾�Cj>;%ؿO����=z��>�p��M$��n����t���ؽ�^�>Un1>c��>�����&>���c��Ϯ�6��>/�t��ܸ=Z��=Z�]>������>��>�[�?����� >{[>��ݾ�J[�������>��r���>=ڎ>*q�>����l�>�>=��W>ф�>�uw�GkW>{�?�޾��/�w�?(鼮�5��_>�ȿ��>��׾�u]<U�(��>-�
>���+���<�>���>	Q�?�=^��?
�%>���b�̒�=�F}>�qx�w�-��U>c~>>���?��=��g>�ɗ����>�3V��Mg>��|>֤�?�QL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       W                                            L       idiL       left_children[$l#L       W               	      ����                     ����������������         !   #   %   '   )   +   -   /   1   3   5����   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U��������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       WCh�@��A���>�� @Ng@ATet@�P    ?���>L/ ?�pA��@�/�@���?���                ?���?T�*@�^�@��(@�@�?�V'@�~?��>�� ?7�\?G,�?:��    ?���@c�@y��@%��?�`�?�V~@?� �?�b�>L&�@{�*?���?B��?�r�?u�=8�                                                                                                                                                         L       parents[$l#L       W���                                                     	   	   
   
                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0L       right_children[$l#L       W               
      ����                     ����������������          "   $   &   (   *   ,   .   0   2   4   6����   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V��������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       W���<��P>���@-F����?�C�>٢F�!)_���4?������P>:�@��\�9RE1�+~=�m����8G?7�޾���u�5?�	��v�#�x@2xu?���UBn�+���Z������'���Y;?+�8���i��An?���?Q�>uW�@�@i-=�eH�Zޜ�0ľ��ƾ�	?9���Ϝ>�쨾�P�2)>I�K�і����m=�yW�$&�=޿Ͻ�&p;�I��,��=P�>�r�M遽�I#=�hJ=$ȩ>�:<���>&��>
g@��C��|�<���>wH���轭2�=�~�=�o>!��<���>x����=�
h��\�=�b> �>#��L       split_indices[$l#L       W                                                                                                                                                                                                                                                                                                                        L       
split_type[$U#L       W                                                                                       L       sum_hessian[$d#L       WD��^CЮD�n�C��BB��VD$��C��C��@��kA��B9�MC��C�H CX�CxS�@�a�?�)A�?���Bn�AD�\C�
CMCn�C+!eA̼�C?$�BIm�CE�A�"9@���A+0 ?���B<�[B�HfC'�,B�B�pB�`�Ba�~B�iA��@W4�B�]FB���B-}#@߅lA�<C<�6A�8A�J�?⋊@�K�?��AL�B7֝?���B��Bd��B��B�ߦA��:@�8B��@?�tB���A[XuB1m2AA.Bٞ�@��^A_�&A�	?��y?��6A��B�oBQBJ�z@�?BuC@M�>@q8�?�X.A6A��C!lcL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       87L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       a<i�Q>=,�P?�>���������k�>�x��&}x<ga׾�l�=CݾƘ��>徽@(>�~6���нI���=�2K��-��l޾��=�q�^Դ�����
9+��t:����>��I>�Pd=w����=����¿�
�A>��;=71>�I���-��]�>S^��I��T">*�r����վ�r�j'���
?�𾉴>U�2���u?	����>�㼽�s�>VU}���IP��K�v��>���>��Ǹ�?6>w����[?1�>��߾�oZ�ݼ�ZӾ� ?����?�I��_y�^þzu9>m1��RV� ὃ�a��>H�
H?�n5���=�n�?>�H=�+���A߾&P��~L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       a                                                 L       idiL       left_children[$l#L       a               	                        ����            !   #   %   '   )   +   -   /   1����   3   5   7   9   ;   =   ?��������   A   C   E����   G   I   K   M   O   Q   S   U   W   Y����   [   ]����   _������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       aBk�TA�d�A���A�`@���AU��?l��A]�@W�&@��C?�� AfG?���    ?�
�A �@�v@S�?8bh@
܆?��,?�:�=�t @�/�@ n�?���    @*?*� @�� @r/(@�?UL�@�P        ?�5?,d�@��    >)` >���@%-?��`>�@��O?�"�@`)7?���?�{V    >�_�?���    >�/                                                                                                                                                                         L       parents[$l#L       a���                                                           	   	   
   
                                                                                                                             !   !   $   $   %   %   &   &   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   3   3   4   4   6   6L       right_children[$l#L       a               
                        ����             "   $   &   (   *   ,   .   0   2����   4   6   8   :   <   >   @��������   B   D   F����   H   J   L   N   P   R   T   V   X   Z����   \   ^����   `������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       a�5n?K�׼^vܾd�>�� ?=Ǿݑ�?�2 ?��|?za��Sw�0��?�*r�����ҿP�=�?]�?U�v�o��C!��\W2�H�J?0ܸ>�i?�ܾ%�4���'�<lgA@^e?y.��8��A(��$>��#�@�'=�Խ�6=���?��?U#�?������ֹ�U�����-?�;R=�r_>J�|�#�@�o�^>�8�=�(�uv>%:}�.�==���d=����� ��q��#�N���=���=üK��~>,�A=.�����>U���5�r����h��������> �U�iK>5%��?^����FV=�P��|hS������u�#�:=p}�%�L�2ھ��=V>d�$<�gk���G�Q�wL       split_indices[$l#L       a                                                                                                                                                                                                                                                                                                                                                           L       
split_type[$U#L       a                                                                                                 L       sum_hessian[$d#L       aD�=�D^\D.�D41C(�$C�5YCD`D�IBў2B�)�B�.�C��~B��nB�/B���D,�B]B�CTA�kyB��A�vgA���B7��ClxhC�B�ϭB1��A��fB�y^C�W�C�ZB�7Ax�.B���A-R�A���@�fcA��Br!�?�>~A�A�AE ?A��Bu@CQ4�A�>B�m�A�>]B~AmA���@s0�A��L?�Y�B�s�Ct7�A��+C�N�A�&!A���A3��@�5A��A��B�}@�%@���A3%�@�gBciC@k�9@��A^�tA |}?�4�@�Us@��
@��?���A ��A�!A�`�C5�A,�:A�� B���A�n�@L�A�T�BA��Aqv?��M@�@��A,2U@���B��L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       97L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       e��ݓ>��,��L> \�>�Bv���!=�L��^�>���>YG�?
��$:���j>�T��<���=�"�>�d>�w����->���?
� >A�[��#��>=��=������.7>�tP� ˌ�KⱽMH�"m��%>_��;���>��M�/`?��>�b����>�R=��I��7����>������n>?�¿�M�ӟE>=W;qo>'��>��Ŀ���L;>P����p�>�PW�dG�>Ộ=�W/?�+��xi>�ѐ>�K꾧�T�/�{>��)?���<��=��r>�[����> ��=d��?���n�>�3󾒩��x>T��1<6�?�o>_m|���Ͽ>�S>�9+��/Ѿ(!�?R\о�,�>��c?[��>�z��_1�?,Q��^gL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       e                                                   L       idiL       left_children[$l#L       e               	                                    !   #   %   '   )��������   +   -   /   1   3   5����   7   9����   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W����   Y   [   ]   _   a��������   c��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       eB�)�A}�`A��A+�v@3~�A�@�6�@�_,@pC�?���<L  ?���@�b�@��L>Ђp?z��?��/@U9!?��?8 �>�4        ?c>�@L�@0��?Н�@K��@�L<    ?|�f?���    ?�?�&f@f�?~�`@3Ɗ>�| <�1�?���>��?7;V=x� @74�?�?vՎ@!�    ?dM ?�]�?�u|@���@�`        ?���                                                                                                                                                                                L       parents[$l#L       e���                                                           	   	   
   
                                                                                                               !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   1   1   2   2   3   3   4   4   5   5   8   8L       right_children[$l#L       e               
                                     "   $   &   (   *��������   ,   .   0   2   4   6����   8   :����   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X����   Z   \   ^   `   b��������   d��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       e�d��d�>L ����y�< �?���??�ȿ�r�.$�>��6=�>�8�>�3_�0�H?�]׿W���2h�>�UϿd�V��+Z�;f�>&��=htn>������?g��@�?���?��P���?��>Y~R�\�?���<lgA?_xI��y���:2@A��i�Ͼ��h�m��ȿ�%��ְM��>ÿ)2���#�ÿ�@;�?�%>��\@D��O��-�?����>ch����>p�<��>-��ò=��G>-���e�R��>��>!�d�b4)<�~�=����6Q=p<�T�>^𽮅%=�$���¾ )�=���P�;[�>7d=�~����=��=�wξ��I�C>|oa��O=�v>n��8=�,�����>Nǹ�Ǥ|L       split_indices[$l#L       e                                                                                                                                                                                                                                                                                                                                                                          L       
split_type[$U#L       e                                                                                                     L       sum_hessian[$d#L       eD�(VC�H@D!��C�lCVs�C�aMCE�BǨ�C HrB0�C6'{C���B���C+�A�d�B�vBqR!B�w�B�+AF�iA�1C4��?��C�vA�mB:�cB0��B�+�B��?A�icA��@���B	�]A��LB��Bi��B��@߶Bt;�@@�{Ak
Ag��@�UC�d.B�G�@�>�AL:�B&A@���BQ}@��@B`YB#�4B���@��l@�H<@IJx@8��@�A�j@d2XA̿�A!��B9��AA'�Bmm?�M!@%wN@��pBn��?��?�G�?�Sb@N/�@ž?@EM:A6��@�@Q��@��^C�٩@�&�Bt��@y�u@��?�^�A/�@p�%B5%?��Bm@[?��Bz@�&�A�%�A�ȷB�}�@��@?ª�?��YL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       101L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       S;������g>!���g�m�!D%>X�R�?��x�!��/�������2==�ި=�7>�����ڕ>�9�^�>��w�j�>_p��͡l>.h>;����~����>O��>U8�>݌c��e=�fT���R>���� R�4� >���R5�3�.>��#���������>�'>��;f��=��X>�t�>���? $��I���>�p�,��?��rிD�>�B�� N>���(��?2�Ծ�>��U>�Te={��Q>��羀�=�na>��	����($>��[�Y 2>�U3���?��>�^�����yO�>��s?dk=�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       S                                          L       idiL       left_children[$l#L       S               	      ����                     ����������������         !   #   %   '   )   +   -   /   1   3����   5   7   9   ;����   =   ?����   A   C   E   G   I   K   M   O   Q����������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       SB��	@�a A��>� @"�3A��AJ&|    ?y�X>��p?p3,@F�@M�@Ȧ�@���                ?��t?_�?ۛ?��G@ w�>�� @��9@{�x@Q�@��?Ub?5o�    ?���?�؀@{?��    ?���?��:    ?�7@���@0�@��@�N@(�?�@E��?�@                                                                                                                                        L       parents[$l#L       S���                                                     	   	   
   
                                                                                                           !   !   "   "   #   #   %   %   &   &   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0L       right_children[$l#L       S               
      ����                     ����������������          "   $   &   (   *   ,   .   0   2   4����   6   8   :   <����   >   @����   B   D   F   H   J   L   N   P   R����������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       S���<��P�,�@-F����?I��>ϛھ�־��4��jt����?�"{?��a�J���<�$��=�x����&���>�� �֢V>�ΐ>�೿(�?�cX@$4>L �>�p7>�{X?2�ʾ�,��ʏ�?�h?�>���#�5��/s?Υ�?�3"�C�;��v?v���x ����?��J?��ǿ��%�@Q!���$q���=��ӽO"K>3�޽���#��=���΍+=��ѽJ}\>Vg̽Ѷ;=��g> �
<�+���a9=�e⽚��<�>&��	VżI��=�Y���F�>��=|>�?=��a��D录�=ޚ$>x�=66L       split_indices[$l#L       S                                                                                                                                                                                                                                                                                                      L       
split_type[$U#L       S                                                                                   L       sum_hessian[$d#L       SD��C��~D~4C��B��Cl�DYSC�q�@Ϙ�A�g�B.��B��Bw��C�
xC�(/@���?��/?�y�A�0 B��@��'B��G@�uB_�@ǿ�CQC�}uC��CkX�A��A\��?�GV@�QBX��Aɹa@��@��A9�2B0��@J�"@D��C2vA��tCU;�B�}�B�[�B��HB�lCћA�CX@�g@��@�UJ@�p�?�q�BSG
?�Z�A�T�@ő�?�`G@Q��A-�@�"A�jA�h?�[Y?�ġB�`�B��A��N@O�.A�ޅC?�-B��S@�xyBk$A�B�@���A�LB�P"C�Q@{҅L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       83L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       _<u�>&�2>�>��=��s���Z�ڻ�>�N>",=�A����??D��
>�3����3>�J�<e�>u�¾�&u>��Զe���=�/=������ﾛa����ݯ�ե�?�����>�qI����>Ĵ��w�h<���)�D(>0�d>�߾�u�=�|B��+�?�W����=�1��	��K-"������W�>��F>�X	�r">N�<�ܓ|?�ƽK��=�/?�q�����>޿��x�r=y߾�0=��-�>�0�#����	�J����V>���<�$=��T����<�Ԫ�҈g<g1�>�B�x:>-�о���>E�9�~Å���Ͽ�=ۆ�����=���?#��=�y�ݚ׽�����CL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       _                                                L       idiL       left_children[$l#L       _               	                        ����            !   #   %   '   )   +   -   /   1����   3   5   7����   9   ;   =   ?   A   C   E   G����   I����   K����   M   O   Q   S   U   W����   Y   [����   ]����������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       _Bp�AkɜAZ1<@�`�A ^ZA)��?��P@=��@J�4@���?�j�@��?s��    ?�� @�@��@6"B>��@�
j?�y�>대?��@ũ5@q.�?���    ?��m?��>�     >�� >��$?���?\�c?E��=���?�:GA�P    >�    >��     >$'�@���?��@�/?P4�?o\X    >^0?��t    >�v`                                                                                                                                                                L       parents[$l#L       _���                                                           	   	   
   
                                                                                                                       !   !   "   "   #   #   $   $   %   %   &   &   (   (   *   *   ,   ,   -   -   .   .   /   /   0   0   1   1   3   3   4   4   6   6L       right_children[$l#L       _               
                        ����             "   $   &   (   *   ,   .   0   2����   4   6   8����   :   <   >   @   B   D   F   H����   J����   L����   N   P   R   T   V   X����   Z   \����   ^����������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       _�5n�a>�^vܾ���?NdL?p]Ǿݑ�<lgA?���@�Z?��*=��D?�ƾq:����@ �ؿ`VW�� g<�i����o��R�0���?��z>v�,?��#8����'�?3�*�� �����3*?��x?��\�p
|��5޾d�>w�=ɼ?�[�7<���7��>'�6��S	@$��g��t��>�V��w>L��o�^>�8�=w�|�uv>뻼to�<��9>?㻽(��+v>�a��Vx<#�r������>�P�Dj �Br�s	#�
g=��2;1{�<*�:�!28�r�;��3����;��d=;�� )�=PƔ�{�=m,���۷�KI��O=�)���<��>DI�=vI������8�L       split_indices[$l#L       _                                                                                                                                                                                                                                                                                                                                                     L       
split_type[$U#L       _                                                                                               L       sum_hessian[$d#L       _D�kgDE@D��Cq�MD�5C䕚C/�C'�,B��AC���BFC��~B��nB�2�B�-Cp AX@�B�/YAwCC�u�A��)A�ߜ@�#�C��B���BWdB��A��OBv�hC�?�(@Ě�@���B,\�A��@��@�+DBM��C׿@
HEAę ?���A�v@	��@p��C�GVA���B4��B8�BRC�?��@mAk�>?���Br|�C��?��:@3{�@U��@���@6��B �'@<�SA���@J%;?��T?�8�?��@�dB	v�A�}�C|�C3vI?��A�οA�1t?�I�@+d�?��uCr1!Aeس?���A��FA���A�1�@޸B	�@�9uBA��?�j�@L@��Aj�@�4�B^6>L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       95L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       W��_�>�;��\�ֽ�da>�P~��3=�c���,�= ��>vU0?�����GF,>GžͶ�����>��j> �`>�j>�5??�X��aǽ�b�������^g=��>�'��M}�1������>e�����>��>���1-��6>�?v=�`�� �⾈Vk?���!<�>�&}=����|V>�����9�>DA?%t>O�ž�'��G��>ړ1�C'>즕����>��W=��
>�c?���>EE���2N<�-��\3=�����u?E�`>";|����=�&>�qJ��⪾I��>������=��4>	��>��C=�#>�=��6?;vʽ��s?�]��>DL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       W                                            L       idiL       left_children[$l#L       W               	      ����                        ����      !   #����   %   '   )   +   -   /����   1   3   5   7   9   ;   =������������   ?   A   C   E   G   I   K   M   O   Q   S   U����������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       WBq(�A��A�n@��@���@�x�@�    ?i�@b�h>v% @J @؋@�Q!>��?�2�    @L}�?��?٫    ?s @��@��?eI @���?�#L    ?_2N?�}�?S��@~j�?�a?T��>�T�            >�) ?��=��p@/�?�dt>�%h?KM�@ R�@]�?�m�?�9?o�A                                                                                                                                                    L       parents[$l#L       W���                                                     	   	   
   
                                                                                                                       !   !   "   "   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1L       right_children[$l#L       W               
      ����                        ����       "   $����   &   (   *   ,   .   0����   2   4   6   8   :   <   >������������   @   B   D   F   H   J   L   N   P   R   T   V����������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       W�]���W��>��.�� g�d��� ??�Ⱦ�?��\>:�f�< ƺ%Ʉ>mf#?��N?��[&>Fڿ �*>�,z�L�>"�j�O�l?y�s�JA� �~>fw�?�$����?*t?'~��o}�>΀�ZR�#T���b�	�!>��=
Ӂ�V��`g@!(�?�QV����a�Y@�}?���?���>��N>��.?aP��V�o�>%�j.�>������=��6=Ƞ>��>�V�;�=l�ս�	+;�7(�;q<�P���z>mBt=B�ɽ�j�=
��>�`�!��qҮ=��L{<�?=%$�>')����<�Q^=��B�>`���>1�p��J�L       split_indices[$l#L       W                                                                                                                                                                                                                                                                                                                         L       
split_type[$U#L       W                                                                                       L       sum_hessian[$d#L       WDq@�C���D��BNFqC�C�i�CHt�A"�B%��C`C	�Cv-;C,��C2�A���B�8@J��B���B_�KA�Ck?Cf�XAt^;B͐iB��,C9�B��AoU�@�A�5�A7�B78|BZWBBQ�@e3k@��@�� ?��CeߔAL�@!�B��2A���@>��B��wB�L$B�'`A�b�A��^@@�x@�&aA�1]@ !�@��@�GhA��A��A�5�A�x�BKQ�?�p�?�r�@z?�o#Cdt�@�T�@���?�g?�HBRB�A��)A��:@�?���?��yB�B/@h�B($�A��
Bj�B�:Ac�d@4�A��<@)
?�/[?���L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       87L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       ];�"R���>1r���^����x>7j��������E>%>�5\���=��=�M�>� ��1�D�׷@>W����>4"�>�K�r>������1>$nS��̫�:_> �=�+�>����>�&Ѿ��<v�m>��G����>?�1��u�>��!�k,����$���׾��>��>��s�X�޿��������U>��=��9>�it=B�>�L�>��>�ᓿ�m�f5?%�����>Ȓ��T����<��ڔ&?�*��u>�:�>�3��pm.��cG>����Ր=0�뾸LV>����1�>� ��i0>���'��>	��m۲>�Ѿ�>P{�?�}>��f��W�>�V%>��J>��iL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       ]                                               L       idiL       left_children[$l#L       ]               	                              ����      !   #   %   '��������   )   +   -   /   1   3   5   7��������   9   ;������������   =��������   ?   A   C   E   G   I����   K   M   O   Q   S   U   W   Y   [������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       ]B�@$��AT �?� ?r��@�,FAn�>�9�?�;P?/G�>+�@	G�?ީ�@�x�@��    ?�V=?���?q�i>�&�?�        ?	��?�?���>�L�@���@#
�@�@)�        =J&�?���            >�        >��?�h}?��?�l?�H�?���    >��/@9:�@��@Q��@<
�@0�)=v��@>��?Q�`                                                                                                                                                L       parents[$l#L       ]���                                                           	   	   
   
                                                                                                         !   !   "   "   &   &   )   )   *   *   +   +   ,   ,   -   -   .   .   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8L       right_children[$l#L       ]               
                              ����       "   $   &   (��������   *   ,   .   0   2   4   6   8��������   :   <������������   >��������   @   B   D   F   H   J����   L   N   P   R   T   V   X   Z   \������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       ]����>�� �,�>��l?:�C?E�v>3u�@-F�?2��>�Op���P>�%>?��a��R�,v������4?ׇa?�@^�S�@@o�>-��/�K?��Ŀ�?���?�cX?R��?�x?�	>��о?�>K>���?@1�>O+����=f1տ��>G���?Հ��~�I?�0��j��f{ۿ'�2<7��v@@r�Q^��G?��D>�� ?�,�g��H4��
���>Fi���=9�|�2ľQt;-�Ѿ%�>?�̾�Z=�y�=�
н�A���C�=ր;3�<S���(h=��v��E=������=����Iw�=$�h���>��3�	=z.>.��=��{�4�=�g`=�'�>	sL       split_indices[$l#L       ]                                                                                                                                                                                                                                                                                                                                            L       
split_type[$U#L       ]                                                                                             L       sum_hessian[$d#L       ]D���Cz��Dn��CjycA���C	DK]�CG�BB��AU�>@F�&B��Bta�C�t�C�F�CBN�@��yA���@�8�A#a�@I>�@Ţ?��B\��A�!B^@��%B��C��1B�Z�C���@���?�1A�+p@���@��?��?�TA ,?�D?���BL+�@�/PA+�pA`��B
�3A�I�@3��@1�hB@]�A犲C���Br�	B�;�A8�CC	��A�R@@6ɂ?���@L�=?�i2A�BGP�?�ZS@C�b?�J~A��?���A��@���@4a�A�H4@[TA�n?�5/?�բB1�{@j�@�@�A�zsB*��Cn{�A��B'�B2JBEE9@���@n�@�[gCyDA��B�aL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       93L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       U<���=��þ�4E>�S���L���\��+ƽV^|>�%�<�����:�����>Vp���t����=�*���>�ұ��u=Q�ƾݹ�<X����Vq���Ǿ��>�3���[�Q�W��>�u��Q�>�`�Z�>��Y���{=������U>B����O�tCC� |��Ĥ>L��?ۿ>�����X>�\>�-��C�>�R��n�>�x����u>���=�1�>��_����?
tL���=R]���=�Ȩ��z��犾>��>�{-���&�#ݿ¼�Ae��7�°��2�?� ��s�Hj>��2�����Z�~?&ƾ]�S��4?�վm�տ��L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       U                                           L       idiL       left_children[$l#L       U               	                        ����      ����      !   #   %����   '   )����   +����   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G����   I����   K   M   O   Q   S������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       UA�4A�*0@ ?@���A�~�?��k?Y�@@��5@��H@��l>� ?9�?�E�    ?�}�@  �    @���?��@�J?���    >ָ�?:    >g�P    ?�@ Ǽ?� �?��`@�@� ?�9�?���@��[?���?�>Y� ?�d>��     ?��l    >fd�>k ?���>�~(>r:                                                                                                                                                 L       parents[$l#L       U���                                                           	   	   
   
                                                                                                           !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   *   *   ,   ,   -   -   .   .   /   /   0   0L       right_children[$l#L       U               
                        ����      ����       "   $   &����   (   *����   ,����   .   0   2   4   6   8   :   <   >   @   B   D   F   H����   J����   L   N   P   R   T������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       U>]R�-�����Rʶ?�b�����QB����?���@�Z�8M�Vs�=�p�!�򾗔n���h���?�b�\�{?p]Ǿ�n;��Z��%ڿ����?�Y����?b]l��rW>s4�o}�>�h'��`g@k��U�r@�>�S޿I���\�X@ 0�@S��腒�Y�>2�L?b]l����<�(���޿3��>�q�Q�=����6�>�E<�m=����k>&%(�)�<|׾ B�=����",���d�[> ���%a� �־j黛F���ԽQ�>8� �ޡ�-#�=�I	���"�> �T���2�q>*Qͽ����"eL       split_indices[$l#L       U                                                                                                                                                                                                                                                                                                                   L       
split_type[$U#L       U                                                                                     L       sum_hessian[$d#L       UD���D�ϢC��C���DC��A�L�B�B�B`5C���D0��B�w�AaܔA
��B�-BtJ�B$�VAnb�Cv�ZAŜ�D(�JA�u�?�r�B��@�
�A	�@�\�@ 9,Ad�B;G�A�� A���C_ЦA���@�I�A�
~D
ZB:	@16A�O+AFaB�I?��l@j,@w��@��@�I @��n@5�B/��A��@��@��"AP7�CP�Ao�A$�AF�2@פ@T��@���A)!D�BF�[A�DZA�ٸ?��B?���@ǭA�V5@�Yo@�3RBysN@)t8@�7?���?�[�?�n(@�D�?�{@��N@)�@?�z�?�dW@�dBhL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       85L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       e��/�>`���t�5=��6>�zb�� �=D�@�l">��	=Ո�?׾��x��"�=����R�>𜾗�>>B,?��.x)>���?o@��·��r)�NwʾK
6>�Y̽�̱>�����r�b�>4*�>M���2�>fe=��>�8�?va>(�=������3=���>�&>��3?����d�=ǭo��D��
#�v\�ر�>�򭾩�.��'=���>6�(?#��>k���:=ʁX?	OT���E�kC��`�>hߟ�8A\?�|>��"�B�>�A����!>"���{�/��$���>����1";>�.[��(��n��F6�>��྘U�>t儾|5���G?0օ>Rn� ��?/wt���(�G�����>�d��'�]>k{K��,�?6��>��?7��j�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       e                                                   L       idiL       left_children[$l#L       e               	                                    !   #   %   '   )   +����   -   /   1   3   5   7����   9   ;   =   ?   A   C   E��������   G   I   K����   M����   O   Q   S����   U   W   Y����   [   ]   _   a   c����������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       eB/|GAF��A�ɍ@�@e��@� @w��@�m�@?H^�>�5�?ѻ`?��@���>���@-&?�_�?�P=��?V
@>��t=��     ?�* ?�?b?�N�?uUi@�}@,T    ?P P@R?`�?���?f�|?ݴ�?��        >��H=�*?#r?    ?h�    ?fB@?
�\?��    ?��F?<��?Z�X    ?��?�h�@
2I>�s ?hB�                                                                                                                                                                            L       parents[$l#L       e���                                                           	   	   
   
                                                                                                                             !   !   "   "   #   #   $   $   '   '   (   (   )   )   +   +   -   -   .   .   /   /   1   1   2   2   3   3   5   5   6   6   7   7   8   8   9   9L       right_children[$l#L       e               
                                     "   $   &   (   *   ,����   .   0   2   4   6   8����   :   <   >   @   B   D   F��������   H   J   L����   N����   P   R   T����   V   X   Z����   \   ^   `   b   d����������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       e��B��d�>��.�z��?��?��??�ȿ�JH��@7>�8�?�?��@=�B��0�H?�Z��<lgA?*�ȿC�NL!�W�������@�}�e� �Čx@-SL?���@ޫ��x?�tN?L�к�a�?�F\���t�C!�?N�>#�B=I���;��iՂ����>α�3�r>"�^@'�?
C��`g�l|�*'Ծ�̦?�=�����=+�?�@^?���?���?2�ɽ�x�<��>$Ř��1���(Ž�@�=��`�]<>�/=��ýi�t>�齟[=Ct��P�:�_��B=���T�{>�7��X���m�c=��ڽ��?=����S�S�>T4�=6�Q��_>R�Y���ʻo�o�=���Is�=�I���5�>[
c=2a�>9ҽ��L       split_indices[$l#L       e                                                                                                                                                                                                                                                                                                                                                                          L       
split_type[$U#L       e                                                                                                     L       sum_hessian[$d#L       eDQ�fC�"C��Ck
�C�C�ԬC{�C�6B�,�A�F�B��vC{�B2vZCDlA���B�9TB��BaluA���Auq�A/�B�?�XC_��A��VBoA@�8�BlVB�]�A>Y@��mB��1@�fBvJ�@���B�bA��&Aݕ@.�AO&|@-�@�^@��*@���B鈇C\�@5e�A��A��A�rNAV�g@��,?��A�A��B��yA4�@3��@`W	B���AN%?�;�?���Bj��@8|;@& �@KQA�EIA��{A�@�@4�MA&�D@ ��?��<?�w�@9&@g��@x��?��ECP�,AC/4?��?���AW^A��A�j�?�y�?��A>r@�Jc?�&ARUAsh�A��AW�!B�N|@��A��?���?��?�*�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       101L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       S;�d��N
=�������==_�>��'��Ѿ���K�R>���S�$=�S>X�>�Q
����%������=�鹾�D�=|C2�����|ZS<��>_�;4\>��=�}j>�En��z>�%Ѿ��}>>M?�ᾠ�d>_d��}�>h���d`���g�wvF��P><3`��F�=�H�>)��>ꦻ�_ef>�/>U@�? "��U��û5����>��(�����v��q;��>���$I����?�*����=��`�8��>�&A��*���>�c=�<!�:��>w�{?�w9��ݾ��>�t���>ѕ->��G��'�>^.�?�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       S                                          L       idiL       left_children[$l#L       S               	               ����            ����         !   #   %   '   )   +   -   /   1����������������   3   5����   7����   9   ;��������   =   ?   A   C   E   G   I   K   M   O   Q��������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       SBNTH@
E�A'-?� ?���@�p�@J!H>�~ ?�:�>��    @���@��@&�x>@�     ?d@�?à?�EO?�>��/?i��?�o@�+g@4�@:G?��d                =� >c��    >h�    >r�p>�DZ        ?�i;@�m?�
�?���@S��@%?�?�L`@&�?��R?�3�>z�                                                                                                                                L       parents[$l#L       S���                                                           	   	                                                                                                           "   "   $   $   %   %   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2L       right_children[$l#L       S               
               ����            ����          "   $   &   (   *   ,   .   0   2����������������   4   6����   8����   :   <��������   >   @   B   D   F   H   J   L   N   P   R��������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       S����>�� ?�VF>��l?:�C�ǮO��@-F�?ӫ�>G�V=��K?l�>�B���Ŀ4�9����4?\�8?@1¿P�,@o�?��@�u�a���?��>r��H4�<���>\ܽ���=��?��x�JԔ>3���2�=�	[>�^�������(�I�ݑ���P"�B�ekǿ#cx�,v�?�@%�v�B����v�/倾����৽�=��d�D1��p���:!�V>��E%���6>'y̾�u<��ڽ]�8=��O��e��'�ӽd�=WG�_�=���>'��8ֱ
���=�$׽?��=��=��"��c=�O_>(L       split_indices[$l#L       S                                                                                                                                                                                                                                                                                                            L       
split_type[$U#L       S                                                                                   L       sum_hessian[$d#L       SD��`CG�,D]��C:VYAZ.D0ڽC38�C�QA�=A0��@%�B���DJaBՔ�B���Cn�@��6AÛ�@��P@䵏@x˂B�&BU0�C�O�Cf��BM�B��?�$B��O@S�?�{�A���@(�?���@;��?�ć@Ąn@%|�?��LBb@���BT�A��wB��C�S�C>�zB)�A��A��IB'�AԈA���?���?�Ou?�,?��?�@�g�?�r�?�x?��@@C
�?�N�AG0.A��@���AU�B)�A�81B"��C��Be�yC�B�@��A�@��@��*AO�|B1@��@�c�A�/2L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       83L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       [<��=�k㾿!�>��7���'��ٖ?>���=0�ν�"���@F����>7���)���/<��~>���=��'���k>~��,���ݿ�H����>ɍ���T��]Am���>���Ε`>�ÿ=Ʒ�=�A辆�?���;�a��a�>Áp��� ����>}����n�>"�𾵅�>���=�����T>e�X>�P^��>�Q���(<����~>�	쾉�o>"���H	>�����=��پ� �����Tj>o������=^P�I�?*��Ӿ��=���=h���	����?����i�>u&����?�==N��?c���(<�C�>�N�R��'��?�u�b���XL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       [                                              L       idi L       left_children[$l#L       [               	                        ����            !   #   %   '   )����   +����   -����   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O����   Q����   S   U   W   Y����������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       [A���Ay�?١�A7�6@�Qx?�v�?Mr�@�eH@��^@|ͺ>�@?$�
?��v    ?�� @�J@�3�@��V? �@@	��@;��?�c�    >�    >1@    ?�D?�C�?b��?���?��@��@rp�?���?-r�>��i?�X?�p@�f�@+?��>�U@?��    >F;�    >x�?cs�>���>fB@                                                                                                                                                                L       parents[$l#L       [���                                                           	   	   
   
                                                                                                                 !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   -   -   /   /   0   0   1   1   2   2L       right_children[$l#L       [               
                        ����             "   $   &   (   *����   ,����   .����   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P����   R����   T   V   X   Z����������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       [>]R>:	����J�?�������QB�T|�?�;R��x�?�ƿY��=�p�r2���n�:e>��?ܭ�=��a>����j�d>��޾z��Vs�%t>�Ӭ��e�?b]l��rW?'~�>&An@}@ �ؿ-��?�ο�̾?Y���?B?�녿 7ľ�����+?�4N��������Q��<�$����<�(�)��3��>�W���0;:�m�	�>
���MR=CN���='�3�աq=X��΍�����(eL=������)<)�`�0��>(2���5d����<��I<����>��U�>-���r�=*������>J<x1�>4v�R;�=>
b�}�I �>����,���L       split_indices[$l#L       [                                                                                                                                                                                                                                                                                                                                         L       
split_type[$U#L       [                                                                                           L       sum_hessian[$d#L       [D���D�B�j$DJ��CR
�A�LpB�C�\D��C��BH�AA`�A8-BJ��BQ4B?�CX:�DR�A��+Aԃ�CJfA�	�A�t=@���@�v@���@SAPo�B)AF��B�_C!�BY9C��"BhlA�``@,&T@���A��B�7B&�q@tF�A��@{�.?�mh@���?��S@��@�'f@5�B�A5M?���A��@�d~C n�?�s"BG@�aZC�<B�G�@�_!B��@�LA��?�8>?�i@%�R@,�Ap�@�hA��B�/�A1eB�?�wG@!�A�/�?��?��-@�?��V@D,Z@��c?���@��@ �h?�{�?�FK@�:�A�%uL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       91L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       i��7����> ���{��V1>�M��h����#�=������>��=�>>�q��n�>�X�����l�=�e>ʖ��k�JsA?&_��[ ;ӗ+>�C>ؿ-=��W���<��=3^s?%��>��ﾒ�?><��$jM>��B��ҝ��&�o�<&k���ۿ>I_/���J=�����ۚ>��>�!�=>�D�$?�2������/�>NAY�Yw�>������?�f>�3����=N��= $?�U�[? ��=_�J?IN>mX%���!>8�̾��O?o��h>�TQ���9���G��Y�TcF>�6����=^!>ui�e�>�����`->�?���6r�yw�>��?!��>9���+�����>��x��f<��>��(�m>�V=�5_?Lq�?Γ��,s?{���G�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       i                                                     L       idi!L       left_children[$l#L       i               	                              ����      !   #   %   '����   )   +   -   /   1   3   5   7   9����   ;   =   ?   A   C   E   G   I   K��������   M   O   Q����   S   U   W   Y   [   ]   _   a   c   e����   g����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       iA��
AU|�A8X4@ʹ�@)��@���@�&>�u@�l@�?M��?�D�@ $h@?�,@YG    ?�@��?�5�?P��?�@�    >��?���>��@�?�Ū?:��?�B�@Z�?~o�    >N��@Y?�_L>C��>ع*?Y�@Y��?�%�>��8        ?��>��>�k    ?�J/>�� ?��	<bj ?!�?�<?h�t?W5�?���?���    ?��.                                                                                                                                                                                        L       parents[$l#L       i���                                                           	   	   
   
                                                                                                                       !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   +   +   ,   ,   -   -   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   :   :L       right_children[$l#L       i               
                              ����       "   $   &   (����   *   ,   .   0   2   4   6   8   :����   <   >   @   B   D   F   H   J   L��������   N   P   R����   T   V   X   Z   \   ^   `   b   d   f����   h����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       i���5�ˈ<��|�4 @�}�"q�>��x>��2?H�?���@4�^>���>z�\?��[@Ⱦ��T��1�?N�@'�=�W5>GH=���6��Y߿a�?p6@�~�%� >���@,�x=̞S����>�x�B��g�?�)8�Nt���\�4�@�=q�l�Å��|yʾ�X0�_�>�o(v?��?�u�?ޟ*?uw�?f\�y��?���>ud2>��>��H����X�<x<@+I>$j��`�>@��<�O�>�^=�h����=]p��f0>����
^r=�e/���E��+�2Dk�~݈=����T<�G=�?����=�P���>�����𽕮\=��x>B�=_ ���轟B�=�L���z~;�GL>C���uP=7h=S9>uUX>>�~��$>#Ǚ���JL       split_indices[$l#L       i                                                                                                                                                                                                                                                                                                                                                                                       L       
split_type[$U#L       i                                                                                                         L       sum_hessian[$d#L       iD7�kC�'�C�J�B�N�CN(gCy_QC6zAח+B�i'CI��@�Q�B�EVC.��B��B���A�V�@��B��A�.>C(O/B�@N�@UlBt�AZ�C�nA���BMY�A��B��7A��?���@�U�B/�B e$A�q�@M�_C [|@�vEA���A�y\?��f?��rBU�X@�SB@��Z@�xA��>C��A�c�@��B7�@���A���A?$B@�CA�.T@Wf�@�ƙ@:j�?��jA��zAK�:A�zm?���?��6A���?�P�?�x?�CzC��?�/@�j�@�HLAӬA:V@�9:B�0A��O@�B�?�B2@���?�NMAW��@�)>C��?��^AL>7@�|@��
?�8Aи�A�U@$��@@V�A/ޏ@�^�A�@t�B7I@�?�U�A���@�l?�j;L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       105L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       E;� ;���]=�L۾��^�_O��d�S>"#��P� �'��W��j�ྱ1w=k>'�?�7�<��G��d�>��׾C# >.�e�ך�=�����v@>�w=Ļ>u�Ѿ�n�>Տ>��򾼝���MB>�u��d>�a9��]�=Y0��:�p>g��>������7>��c�۟=V��W�}>�T�7]>���>#����>��A���!�
{3�4����
�>�<����e>
��>����6���
j�>'�a�p��<�G>=������=�N�>�i L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       E                                   L       idi"L       left_children[$l#L       E               	            ����            ��������������������            !   #   %   '   )   +   -   /����   1����   3����   5   7   9   ;   =   ?   A   C��������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       EB�'@eh@��">�@?�"�@ӎ�@�2@=H� ?>U    ?F�a@��@ �@�!H                    ?N
?r��?��?$o�@=�?���@Y�@VFT?��?aC?A��    ?_    ?]�    ?c�L?��@�j?�I�?�Ej@�M@��@6��                                                                                                        L       parents[$l#L       E���                                                           
   
                                                                                             !   !   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *L       right_children[$l#L       E               
            ����            ��������������������             "   $   &   (   *   ,   .   0����   2����   4����   6   8   :   <   >   @   B   D��������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       E����>��l>�]9@-F�����U�*@��@V*ʾ��4��!? P�?�s}�%�>���>av�R��Ž�x�=܈6?7��?���@*��>�&�@V۾+�������G�?\�8���ڎ��V����d=�L�@��>#��X���a�?=�`?=���+C�<��2�^R������<��X���> hf�[�=>�b=Dy�6�=�(N���¾&-q�X���s=�{ѽ�M�=&�2=��[Mw�&�=IBu��Tr<��=cg	���<�+�=�J�L       split_indices[$l#L       E                                                                                                                                                                                                                                                    L       
split_type[$U#L       E                                                                     L       sum_hessian[$d#L       EDw�ZC"d�DN�*B��Bv�CuKhD�PB��r@xՎAR)*A���Bj]C:�QD`zB$m`B��G?�
�@+��?�[9An�#A�BH��AJ/B�.B܄tC��Cc~�A6>�@b-@܌�?�)
BC�+?���@�N@,��A��B?LBW$B�X�C8��CFeA�=�CK��A�<@Q2o?хd?��?� �@��?�`EB<O)@��@h*AH�mA��hA���A�o�Amp�A���Bzg�A'A�v�C(m�BF{iB�OAHzdA4tB|wqC�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       69L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       K<l[	=L����/=��A�'f��H�ڨ!>@��(���YB��tm��ǒ=��ƿ �����>v1e=	=<w�o���1>41/� �ھ�%�g�>�����1n>��/�Ǘ�>�]����>��A���y=%����=(������>�]��uؽ�g���~>;!���>� <<�4{>�G��֐u=w)O>�9���<�Ye>�w;��#>m	�Vs<�X	?Ĩ<ɸͿoi>ލ ��˾�wd����>������ѿh1>V�̾�K�=$5�@멿*��O�>����>��������L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       K                                      L       idi#L       left_children[$l#L       K               	                  ����   ����               !   #   %   '����   )��������   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G������������   I������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       KAt��A3��?�@�`�@In?J��>���@gǄ@Eg.@%>��    ?5�@    ?���@sr�@Wb{@A��?L�H?�Ţ@QY?�p�    >T��        ?Ug�@<�x>�Ȭ?��d?��6@k�?��4?X}K=���?���?(�@@��@'b?o��>�V0            >iV                                                                                                                         L       parents[$l#L       K���                                                           	   	   
   
                                                                                                           !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   ,   ,L       right_children[$l#L       K               
                  ����   ����                "   $   &   (����   *��������   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H������������   J������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       K?
�>:u�*�v�/?��I�'�QB>��@	~~�gJH?�ƾ�%��p�n�����?O��Ѩf?L�>�J?q��h}�>��Ik?�ѵ��n�=ہӿ#Gx�T|�?%�?�R>�T=������ٿ; ��h ='�"?fʿ 7Ľ�Zܾ��=?�q�>3X;��=��B�[�<�K�=�=�k<�==��H:���=�8��/��;�?>,��;���)��>��֎��o��D�>�n��qȾ"}=����<D�@�g�2�&�Y��,�>ݾ��=)M����]L       split_indices[$l#L       K                                                                                                                                                                                                                                                                             L       
split_type[$U#L       K                                                                           L       sum_hessian[$d#L       KD��~Dp��B�C"D@�CCj�AOB�9BC���C�9oC
kB%�a@��@��B�#B�`C��BB��C�L%A�ԟA�tB��8A��+A�6�@jH?�n?�"�BHC���A�B�B��rC�`�A��"@a�A���A���@��IB�<B.2@��As��@<;?Ŏ?��B�HBv!dC���@Շ�@$�A�o�A.�A�kB�O�C��V@��O@��A@v�?��X?�8�?���Au/�A�@�Wy@jbJ?�t�A�;�B��-AGpkA¤.?��U@-��Ab��?�
IA7��A�!L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       75L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       g� �Ͼz��>
�ʻѽ���%�>�-����ӟ=ɦ���v�>���=��v>պ���D>�����形��<�}>��J��C��2�$?,̽��A=m��>���>��H>8���m��=5�?M�1=�ǩ�N)���L�>�����*>�ھ1�m>�d��J'��[Q����<g[}���>:���|�=�kܾ���>���=�eZ=I�h>��~���>�SӾ�!F= |�>���c/w?p��=#">c�꾽׼�
���= �>���t5�?x2>Y9�?	M[>ED����>���B4?Eb1����>��3�t�j��::͸�1\>����o�=�餾楹>��? ��=O�i��>�+>��=B���w��	�>�c�y����s>�Y/>�V����>�G2?��L>�V�[#uL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       g                                                    L       idi$L       left_children[$l#L       g               	                                    !   #   %   '   )����   +   -   /   1   3   5   7   9   ;   =������������   ?   A   C   E   G   I   K   M��������   O   Q��������   S   U   W   Y   [   ]   _   a   c����   e����������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       gA��MA)jA�@�՛@Ѐ@��`@���>�{�?�u&?���?!�j@�?��0@-�|@΄<�	 >���?�&�?��D?P#@?�c
    >t�B?�YZ=7 ?#��?���@:/`?��X?Q�x?hy�<��            ?��[?�D�>6��>��?8� @,T?�'s>�1�        ?�Tz?�J        ?F�>�j�>�Sn>d%x?S�h?� �?��?��>��    ?W3                                                                                                                                                                            L       parents[$l#L       g���                                                           	   	   
   
                                                                                                                           #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   -   -   .   .   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   ;   ;L       right_children[$l#L       g               
                                     "   $   &   (   *����   ,   .   0   2   4   6   8   :   <   >������������   @   B   D   F   H   J   L   N��������   P   R��������   T   V   X   Z   \   ^   `   b   d����   f����������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       g��(�ˈ�����4 @�}�;�1@��?F�?H�?��@@4�^?xc���`>��x@,$���?�o����?N�@'�>�q>1�\=����(~>���� hL=���?��>���?"C>9g¿;Y��a=�Gy��� >΀����?�8?�)8�Nt���\�4�@�=_T<�����g>�8�>͍=�j�FY?�0W?
��>�Ӭ?��3>���?n:�>޻X?
X<C��@Y�'���6��ӽ�H4<��=�E����>!]	=�U�>$�:=l����K�=7T��S>l�;��N=܇q���@��¼��*��no=�T�vB<�~ž
co=�ރ>�J<,���e=�f�> h(<i���
H���=���>+����=��=�5��˥>�>�#�=�hA��{�L       split_indices[$l#L       g                                                                                                                                                                                                                                                                                                                                                                                  L       
split_type[$U#L       g                                                                                                       L       sum_hessian[$d#L       gD#�_C��aC�6^B��C.Y�CO��C ��A�>�B��VC**\@��^B�9�B̒CM�A��8A��@I�B�|�A�}C
A�ʓ@ m@i�B��Aj^~B�WWA���B��jB�Д@�aAP��@M	A��%?� �@�QB6[0A�<{Ao��@I,BC�@� ?Aw�wAY�?��t?���B�J@�AY�?�^N@j!VB�L@��AFS�B5�pA�l�BGJ�A���@�W�?�O5A*�c@q?���?�bA�vAi=�A���?��@��uA+�.?�X�?���?���Ci�?��@@��/@��A��A�@��VBX�VA�V}@���?�m�?�,K@0B��@�2@ȑ(?���A"�@b�Bp�A��A.��Aw߮A�`ZA�5a@�6A��@@�@7�A ��@&�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       103L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       M;�B����/=�(����'�H��=P�v>�җ����~x���#�P��-��=�sn��>��ÿN1�M�*q�>�ݾ��0>@|M�X�>o���_�>���=�yp>ԾT��}�>�����>�]:�ä<�츾�G>�6����T=0��=�W>�䆾�׽��y����>�~.>F��>�޾���>(r�B�>�L�>_~�ȇ=���?⃾��+�*8?%Ծ �=	���ڸ=W�?pҾ�)�=��#��L=� >%�x�	,�>#�?˛���<�x�?������?�k�%�j>�a�?&�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       M                                       L       idi%L       left_children[$l#L       M               	         ��������               ��������            !   #   %   '����   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C��������   E   G   I   K��������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       MA���@`@�>�v�?�QC@�h?�d<��         ?	�@3 @~J$?��?B/�        ? �L?C�p?��L?q��@���@"9�=��    ?�&�>�%�?� >���>��=�K@?��h?��>9��?Q�@��@���@bSl?E�        >�8>�n`?W�#>x�                                                                                                                                L       parents[$l#L       M���                                                     
   
                                                                                                                       !   !   "   "   #   #   $   $   %   %   &   &   )   )   *   *   +   +   ,   ,L       right_children[$l#L       M               
         ��������               ��������             "   $   &   (����   *   ,   .   0   2   4   6   8   :   <   >   @   B   D��������   F   H   J   L��������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       M��8\>��l?ܭ�@<������n�\�@R�������j�? P�?�x�����=���>�06�]սu*?7�޾�*?�q^�����#cx@{6@��=�r���_�9�?��p���>k�>� >����?�}澒T)���,@^e>�o[?�^=>��x�ϵ��ƒ?)�n@w\�d	L�4}o����=I�#�h�=���=)�˽�<��1>!ܞ�D�8�w>�̽@A<%}��;7<���>#�����<������f<矚=F�*�$��=DY�>�!�	��;�]�>����>`�G*=�BB>.�L       split_indices[$l#L       M                                                                                                                                                                                                                                                                                 L       
split_type[$U#L       M                                                                             L       sum_hessian[$d#L       MDdp�CN�DC\�B�	pB)D0�B�-Bġc?�XA&QOA�)�B���Di�@�%�B���B�?�j�A]2�A ~Bi��A��C��C��~@6��?�r�A1�1Bw]XA%��@]�&@��2@]]�B*�Ah@+�AZwB&<�ChK�C�=�B='?�Y@?�ʧ@�E�@�̠Ad�BO�A
�a?��Y?�&?�.%@'��?��?���@��A�1Al	+@{iA@��?��1?�,�@�s @�z�A�$�A"�^A�r�CL=�C���B:
oA&��A��X@;�?�@�.<?�y�@jԛ@�_�A�_RBuL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       77L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       E<z�x=O�-��"=��s���u�������>�*'=-�i>Y���ψ��w�>�P�8ؾ��d>�5��r7;=�	���,>��`�O����jl�1�:X�ަ�>� !�����:1���u�>�n�>��=��{� ��=é���K��K�����>�P�<����M����>��ԾN�>�kn=_(���-?4�T>�r�+�C>�n���>�Ji�nj���>��=^G���r¾�E�>�h��A�>S�\>�Ѿ�&վ�5�=�uj=�b{?Z�>sվ�?OL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       E                                   L       idi&L       left_children[$l#L       E               	                        ����            !   #   %����   '����   )����   +����   -����   /   1   3����   5   7   9   ;��������   =��������   ?   A����   C��������������������������������������������������������������������������������������������L       loss_changes[$d#L       EA@�A�t?���@�z{@T?'3~?;3�@#��@��C?��>è@>�a?C��    ?K��?�i?g�@��b?y�=��    ?@�p    >���    >�,    @6�    ?��p?��>�j'    @�f�@&�@*�?'�        ?� �        >��=�@�    ?��                                                                                            L       parents[$l#L       E���                                                           	   	   
   
                                                                                             !   !   "   "   #   #   $   $   '   '   *   *   +   +   -   -L       right_children[$l#L       E               
                        ����             "   $   &����   (����   *����   ,����   .����   0   2   4����   6   8   :   <��������   >��������   @   B����   D��������������������������������������������������������������������������������������������L       split_conditions[$d#L       E>]R?�2����c'�h������QB?K�Q@�@/�@,�=�Vs�=�p�D7>�]��� g?%�?|�G?�F�?
��y/�?5Um�+�6<lgA��E�#�&��<�>�a8��"@k��V�^�M�k��	������<�?5�J@V�>
0j<�����?��e=ˁ̿#��L��<���?8�>X��>D��N'=�����P==�&����9�=1�<�^7������S�>mؾZ�=}�=3�Ƚ��g���<���<�v.>!9�= $����_L       split_indices[$l#L       E                                                                                                                                                                                                                                                        L       
split_type[$U#L       E                                                                     L       sum_hessian[$d#L       EDs#�D\�6B�,DN�Be�@A�q�B�O�B�/�D0Y@�m%BM��A��@�A��B"�#B���A�^D%��B,��@���?���B��A_�3@���@�f�@��M?��)A�AP&mB��6BuU@q�@@�D�eB�J�A�,A��\@Y�4?�Q-A�ȠAym�?�{�@E7D@XC^?�2zA�N?��B��&@~B	A���AB�@%o�?���B�t�C��B��BK��A�"@��(A�\�?�˔@�\AA�1�?׋�?���?�Ka@�@�2�A�zL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       69L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       e����l'=�2Ӽ@�'��-}>h ���	��X�=��
��x��8�,>1>��Z�K+
=�N=���˽�|=�a?{̾�(U��0پ_&�>�C����>���>��h=�@���e<��=*8?]> S���D-�5=�>�ڴ=�H:��İ?`w�؍0�ΣC�܂�>�������e/�>��O>�Ҋ?䥾��%>�L����<D,�>#��Q�J��.�>8��?H��'j>b�h���	���b>���>�X�LV���t!>�k����/=�
O=l�����>F$������H�?3�����=��׾�>�z:>�v�=�)�>��㼌�?�>t��=`Nv� ��? ��=-,�=�<���(���m>s!%>�w@���¾�Q�>J,>0V����>�l����P?J!O>�{�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       e                                                   L       idi'L       left_children[$l#L       e               	                              ����      !����   #   %   '����   )   +   -   /   1   3   5   7   9����   ;   =   ?   A��������   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       eA��A5,@�k@n�?���@m�@\%C>�k�?���?KE ?g�@T7G?��(?�;6@��    >�|&?�+    ?Ka�@�?d��    ?뽉?���=���?�$�?$F8?eL�?���?�4=N(z    ?��?�]�?��?4�@        ?L�{? 
�@�|@+d�?8`�?lr@?/��=Y >�w�>S�(?:�?k�?"�B?4�@6n�?�-}>��8                                                                                                                                                                                    L       parents[$l#L       e���                                                           	   	   
   
                                                                                                               !   !   "   "   #   #   $   $   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7L       right_children[$l#L       e               
                              ����       "����   $   &   (����   *   ,   .   0   2   4   6   8   :����   <   >   @   B��������   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       e��(�ˈ<��|�4 ?���:2�>�<>�����p�@'�@"�>~|>�K?��[@Ⱦ[z���?#|>���C԰��,�e� =�궿��ſU`�%[�? �*?��P�%� ?E�?�ڿNt���j?�:[?�K>#�@�}>?@���P>�q��,��o}�ZR>�ʜ�i��"*�<��>�v?ޟ*��|�9.	?U�v?�[�ڸ~?2V�@.���@=����<���>��=���u4㽯��=��7���<�?�<������h=! ����	��>0�=��5<��Ͻ=�_y>	3<�˖>���>$JZ=��"<��z�=�>��<O�"=W7��d��8�=��=��M��x����=�5=S�8�=c=��½�W�>r�_=�-�L       split_indices[$l#L       e                                                                                                                                                                                                                                                                                                                                                                         L       
split_type[$U#L       e                                                                                                     L       sum_hessian[$d#L       eD��C}�nC�1�BϪIC�ICD�C��A�N�B�֊B��B��Cd7B���B���B��Ak��@��kB�:`@�¢B��@΀BfU?�ԚB�W�Bt�+BV�A9��B'�A�R�BwU<A ;|@�V?�2�BjΛA�LG@��B�P�?�Oh@��EAĂ�A@�0A)<Bn`�AP&�B@�zAYY!B �p@�ĭ@��B�@�_rAv��A( A�ǖB�qAOf?�`�?�q�?��B\ @l� A�΀@S�:?��2?�W�B�FR@MLA^eA*�?���A/��@
y;A��A��Bl�A+L�@g�Bw�A�A}u@sn�B�b@?@�@� @0�Y@�j�?���?�^�B?%?ߝC@L�C@�tzA�v@�@L�`A|��AY HA��@bI@���@�� L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       101L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       A;�ށ�ҘN=�����N˾/��=9'>�kѿ �|�0���l��R`����>�Y=b	�>��u����֌��e=�X�k�=M�=��>���>���7�>ux;?����ht��S�?m��Xվ�{��q�Qe"=�s�>^8���<����>����e>Wd�>F\>�~ؾW�>}�,� ����-���0p<h��Ǘ��e�n8�=���>x�1��N{��<���#ȡ>�e�]<�>�s������&>�z�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       A                                 L       idi(L       left_children[$l#L       A               	         ��������               ��������            !   #   %����   '   )����������������   +   -   /   1   3   5   7����   9   ;   =   ?��������������������������������������������������������������������������������������������L       loss_changes[$d#L       AA���@�@�R�>���?�l�@R�P?��<<^�         ?	� @�#�?���?�)j?V;        =���?[n@aj@]S�@vh�?�R(    ?��$?$��                ?j?���?�<?�"�?���@�@'x    ?M�>�[�?x\?�<�                                                                                            L       parents[$l#L       A���                                                     
   
                                                                                               !   !   "   "   #   #   $   $   &   &   '   '   (   (   )   )L       right_children[$l#L       A               
         ��������               ��������             "   $   &����   (   *����������������   ,   .   0   2   4   6   8����   :   <   >   @��������������������������������������������������������������������������������������������L       split_conditions[$d#L       A��8\>��l?ܭ�@<����?0\�T�z@Q��S��Ae�*<�h�@�Z�h88;�A:�l�*4�>���M��>��b?�6Ŀ"*�>���9ND?��P>���q༼�>O�>��?{(b��K����N��@@W��1�N��X���>�Cu������>嵽�X=�#��1����;��D��#�/�z����<� �=�"���*��9�;�ؽD�[>�
�1�=;&�K>�����=�,�L       split_indices[$l#L       A                                                                                                                                                                                                                                          L       
split_type[$U#L       A                                                                 L       sum_hessian[$d#L       ADU9`B��D9��B��~A蹾D)KB���B��P?ȋmA#@A��C�<CN�Agn�BS-�B��?�4@A0A���B�i�C���C3��A�X�@��5A'<Aܞ�Aɼ�?�h?�&�?�+�A��B��B=#B7�*C�TB�Bj?�CoAʄ�@��O@�l(A���@�_Ah�@�v�A���A�QA�B$[A�0�A�w{AH�C���B��.@��IA>bB:�?���A�i@g��?ۢ@w\>?��$A&�
A ��L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       65L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       =<m3,=7L����=��{��5P=��1����=�ҿ�$��>J����Ԯ>�~���L�p"�jt�>*N�bY=��&����>�0�{����<=����$
>A��^�����>vj�=��%�̝���N�C�g?銼����͒�>�Խ�P=P�����]<
�b��?�>��?=~��I=�k����><�I=�;ь�=�w�x�r?+�½:Ӿ�a�>�Tk>{����վ4|þ�$���?#�cL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       =                               L       idi)L       left_children[$l#L       =               	                  ����   ����               !   #����   %������������   '����   )   +   -   /   1   3   5   7������������   9   ;������������������������������������������������������������������������������������L       loss_changes[$d#L       =A-�@�D?�&`@�&�?�O�>�Su?���@���@O^h?��>�2    >˄�    ?��@���@UC?�|�?�>�x�    >�             ?��F    @U�h@4�@8�?>?n6�?Ϡ?�!?���            >�k�?��,                                                                                    L       parents[$l#L       =���                                                           	   	   
   
                                                                                               !   !   "   "   &   &   '   'L       right_children[$l#L       =               
                  ����   ����                "   $����   &������������   (����   *   ,   .   0   2   4   6   8������������   :   <������������������������������������������������������������������������������������L       split_conditions[$d#L       =>]R?�2�Yq`?΄�h�<lgA�QB?^�#v�?�@^@S�=�1��d�����>�6n�&�M���j��N�?
���T�8M=�-���=h�w>�]��8�?v��Q�~?���F|�?��r?]M�V�Կ5ΐ>qL�5�<zgx���\>�)���=ń�<��[�<��=@@�s�=b��=�{��u�=Gp��!�>N"�_P����=�eN=��V�d��X���7|��z�>D�DL       split_indices[$l#L       =                                                                                                                                                                                                                            L       
split_type[$U#L       =                                                             L       sum_hessian[$d#L       =Dc��DP�B��%DCĥBM��@�QB�� D0WFB�j�@���B6��@%b�@V��A�b B(x�D��C*y1B ��B6@�q�?��B1@5?�o�?�:1?�	;A�C�A/\iCh$�C�_�CA�A���A�!0@�A�AU�B�@Q��?�M(?С�B*�&A�9cA�C5�B��BB*C~4�B�A.BH��?�EA�w9A]�A>��@�.�?�M@���@��?�\�BԹ@�cB�A���?��hL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       61L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       _��ʗ�[r@=��;�N��9^>=�&��mҾ�>i≮о�S�<E� =�2x>��^�J=��<�!h���N�:>�a��S�R����?�,��`<���>��>�s=�F�>غ��9�<��v?����5��9��x5>Z�K����>��#� �=}�I>��+��Z=�kܾ�N�>̝�L8>a:O?���@�>��#��e�>ЧѾ��^� �j=�K����<«I��/�>��龨�5�Ҥ�>���>�P�yX}����PP>�
���d�R�¾Ԕ��D��=��۾吳>2�>���?I��qyb>���>ԓ���Ɩ?��=>���%ٺ��T��xS>��ѽ���?%�A�L�1��w��<��>��=�?/Z0��ب>���L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       _                                                L       idi*L       left_children[$l#L       _               	                              ����      !����   #   %����   '   )   +   -   /   1   3   5������������   7   9   ;   =   ?   A����   C   E   G   I   K   M   O   Q   S����   U   W   Y   [   ]����������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       _AY�h@�z@��?@Sl�?�8P@ay�@ �>y̠?��L?_��?\� @U�?�>P?e�l?��f    >)��?��    ?�'?B�     ?%�?�o-?��L>e�?���?���?���?�Bp            ?��?�� ?UFP>��;>�!�=D��    >�B?x�s?�I�>��?Ġ�?/n�>6T =��@??,    ?�>d� ?�י?��?W,�                                                                                                                                                                L       parents[$l#L       _���                                                           	   	   
   
                                                                                                   !   !   "   "   #   #   $   $   %   %   &   &   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   2   2   3   3   4   4   5   5   6   6L       right_children[$l#L       _               
                              ����       "����   $   &����   (   *   ,   .   0   2   4   6������������   8   :   <   >   @   B����   D   F   H   J   L   N   P   R   T����   V   X   Z   \   ^����������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       _���5��n>����&��@ n�?}��>�$޿R���Ѭ¾+��@Ij��4�>ͻտN�@R<G??���?�F>�@�(@�}>)%��.F�w�ʾ{ܿ9�?��h����?�>���>9kO�����V�>��?�>@���/,@N{@=�9�>�3_�o�>?O����?�[޾i�J@I�L?��v>TZn�٭C?O��?U�v?�D>ud2@;¾;�X��Ҟ=��K��R�����=�+�>c���������``=>�s���x�}P����lJ�=�Q�	�9=V�=���>%)���n=�ǘ=������> ��<d�ҽGF�(똼���>O~��cc>F��u�վz��bI�=�Z<8��>Rl:��jd=��ZL       split_indices[$l#L       _                                                                                                                                                                                                                                                                                                                                                      L       
split_type[$U#L       _                                                                                               L       sum_hessian[$d#L       _DA�Cd�C�s�B�B�-�CSp�B��`A�xB��zBÅEAD�CjB`�B2^�BS}�?���A�o�B��$@�EaAz�\B�%Z?�z�AUJB�X�BR��B*�8AV�@�:�BWlBE�0@\��A�O>?��B���A���AO��@,�B���@�@�@̷�B�%�Aa�B`|A�,�@�tB�@bQA�j?�sj@l<A���A��6B")�A(�Bj�NA�S�Ag�R@?��A9'?�M?�j�?�X�?�"�B��Q?���?�c�@"��@v��A4�B���A)J@a-�A�_A���A'�R@� @p:.?�[�B�`?�J�@�1?��?@1Z@ⲧ?�2@��@�sA���AH��@e�0Bq�@��@�=?�)�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       95L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       7;�߮��u=U������D��vN=��S� �^�vx��	Խ��+��.<��=��f>�Ff<�i����5���;>�N�=8�����)�=�WW��8>�澼�>��o�=�\>��<�y}��hԽ6#���=$�->I��ݦ�>�ND��
;�[��X>M�"���?;�>�9��_F�oǽ�Q�>�=��!:����j�$=��u����=o�P>��!L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       7                            L       idi+L       left_children[$l#L       7               	      ������������            ����   ����   ����            !����   #   %����   '   )   +   -   /   1   3   5��������������������������������������������������������������������������������L       loss_changes[$d#L       7A�W�?w�0@z>�<� >�s�@vD]@uݰ            >��E@1�?�+@�    >�W�    ?���    ?곡?-rD?�]�@'�"    >�B�?i3�    @	?͊h?o>�T?���>���@�z?�P�                                                                                L       parents[$l#L       7���                                               
   
                                                                                                           !   !   "   "L       right_children[$l#L       7               
      ������������            ����   ����   ����             "����   $   &����   (   *   ,   .   0   2   4   6��������������������������������������������������������������������������������L       split_conditions[$d#L       7��u@?:0>�]9@M�3�	\ͽU�*@���nq�-Z���@2W@=�D?�D�H�'>���8����@'�>�?�Ù;�l��S�>��޽�v?v�?�C6=�҆>�s��?kª?�r�?KN�?�7z���^��7���>b)� w::�mY�ǜ�=w2)�#��>�=�D{��rT�(�"�dE=�@�ADF�Ϣ�����=	Vz��1�<��0=�J(L       split_indices[$l#L       7                                                                                                                                                                                                   L       
split_type[$U#L       7                                                       L       sum_hessian[$d#L       7DG�B� �D55�Br�LAf.�CX��C���Bn�\?�=�@�LA!�bBQ��C$q3C���A���A��?�n�BFE@9�C��ANɰB�rC�S�?��G@�PBA4�?�
NC �A�O9@�~|A�rA�
 A ��C�{CC+�B@��?�$�B*Y�@���B��BccA%��AP��@Ǻ?�j}@��@�@�ZA�3z@ٕ~?�@C+YrB�:'Bp�'B���L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       55L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       7<a�z= �s����=o����yܾe;Ӿ��=�.��;-�D:o��x꾊Z�>~Y,=Ǹ����<������&���h���~��1
���� �ھ�-?�h>�<�{����F�ť޿v���p��>���>5*���q��Α=:�?+h;>��=�*�>�^>�����>�)���Ծ[�V���>Ц�����։Y��3:���>D����>�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       7                            L       idi,L       left_children[$l#L       7               	   ����                        ����         !��������   #��������   %   '   )   +   -����������������   /   1   3   5������������������������������������������������������������������������L       loss_changes[$d#L       7@��@�2T?k��@k�/?@5P?u��    @C�>�:�?�|�=(��?��l?N2@3��@,ʹ    >o��=Ǯ ?v]�        ?��K        =J]0@��@5ZP?�n�>e�                ?��>��>�R�?���                                                                        L       parents[$l#L       7���                                                     	   	   
   
                                                                                 !   !   "   "   #   #   $   $L       right_children[$l#L       7               
   ����                        ����          "��������   $��������   &   (   *   ,   .����������������   0   2   4   6������������������������������������������������������������������������L       split_conditions[$d#L       7?p]�?g(?��@$> ݼ?�*F�M�?a���3�a�QB?��2>���?s:������*;��x�Xň�e�n=N�h����Ӿ֡��9��Ϸ?䵂����>{Dn�#�x���4�#X���+T���k��-�Vխ?���?��>>M�G=5��<�3=��q=�ȼ��C=(��L���g�b��4�=�a��1�� �ϼ���=l��7L       split_indices[$l#L       7                                                                                                                                                                                                         L       
split_type[$U#L       7                                                       L       sum_hessian[$d#L       7DV�}DG��BnʚD=&4B(I�BzA�v@D9�AdE,A�Al��Bf@J��D�0B��s?��{AL�A,U`A��W?���A\��A���AO�y?�le@ `~C�d�C�W�BҎuA���A-�V?�Z6?�'A�A9*�@�p@A@Aa�?��m?�&�C|.�B�4�B�'aC��B-�BwR�A(AU�@���@�m!?�0@yH@F�@�$�A0��@D��L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       55L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       [���Q�C+I=��k���־ϴ=>!U-��ĺ��u;a����Ez<���=s�K>�����0=�Y���)>��=h�3��$�����>T�
����>�D~;�N�>�&�>���>JS��y�=�����>��W<B�J����< s�>��{��Ľ�Mľ�a�"k$>l��iL?`u�lƂ=v�׾�>�>�~���ν�h(>� `>;現�ľ?)���G����}=�[>���������>��c>�~��HE>D�?e>9�]������KR� �p��v�>]���e_�c�P?�t�eX����>N���=�^�>��վ���>�?ӽ�W���6E���>=|�<�ۿ�>x-��Jo?oA��xL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       [                                              L       idi-L       left_children[$l#L       [               	                                 ����   !   #   %����   '   )   +   -����   /   1   3   5   7   9����   ;   =����   ?   A��������������������   C   E   G   I   K   M   O   Q����   S   U   W   Y��������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       [A)��@��@:��@=��@�@6�8?�Q%?�ZP?�;�?6 ?nz�?��>?��?l`?��?.Gp    ?��D?B$>�+�    ?*^?�X�?��?�:�    ?�?�?ket?���?0(�?aP�>�RI    ?��.<+�     ?F)�>?π                    ?�}�?-��?sC>�g?��?�� >l�J?rH    >��~?O�3?�?? �(                                                                                                                                            L       parents[$l#L       [���                                                           	   	   
   
                                                                                                               !   !   "   "   $   $   %   %   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   4   4   5   5   6   6   7   7L       right_children[$l#L       [               
                                  ����   "   $   &����   (   *   ,   .����   0   2   4   6   8   :����   <   >����   @   B��������������������   D   F   H   J   L   N   P   R����   T   V   X   Z��������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       [�Ke�<�h�>,��@5
�sb?��2@-�>J�y@XT����?�n� i?c��?٨���=�໿.$�?4Kd@;&�=Ps@lb>X=Ҿ�T�?�@^>G�%Ʉ�?�?&*h?�	&>G$��D�6�>qѵ�C����/��B��=������>(s����>~|�%�Ҽ�@`]� }b?��J@4�^����>K�?�
�?b]l@�?9�:�����qt=�V=+
1��#�=*��>F=^�׽��&�-2�6 ��[.=���	�����>(�����7��%�=w6þ6I=�=�{ͽ�U�=�d��K��=RӾ���ȅE=cbQ<��/�=�͂�ȿ�> ��\�L       split_indices[$l#L       [                                                                                                                                                                                                                                                                                                                                   L       
split_type[$U#L       [                                                                                           L       sum_hessian[$d#L       [C�LGC_mIC���C`jB��CT$�BlhA�yB��B�ǆA"��B�_�B��&A���Aڇ�A�  ?��BƎ�A�O�B���?��@�@�sB�m+A��A�%BpǸA�G�@͍AjTAJ��@D��A�k�B��HAzHA
�A�B��@�?��@mT@a)x?���B�_�A`m[A�/�@�i�A�1�B0.�@AA��?�)�@�£@��D@���A511?�S?���?�hBV�BN��?��J@�G~@���@~�@r&B�<Bf��AA��@�w�ANL?@pL.@uQ@��@`}�AJC�B&�b@!?��?��@��ApY�@o�2?�<&@��@w�@�l�?���A�v?���L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       91L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       =;�e���2�=7����F�9�=<� h>��z��f½��!�'`�=2���P9K>�/<�Ts������=��o=��>��ϖ�=�=HP�>��f��>Q�\��*�Uy>w�A�
�=��=T��x(�>ҵ�$>�.e>'�Y>�|���n%��r]>����!��(t
�蕾�!)=��ھ���>�����<�ނ=m5���:�F�S>�C�ކ����>�t����>�HO�@?�>�&�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       =                               L       idi.L       left_children[$l#L       =         ����      	   ����                  ����            ��������   !   #   %   '   )   +   -����   /   1����   3   5   7   9   ;������������������������������������������������������������������������������������������������L       loss_changes[$d#L       =AV$O?f4 @T�\    >�{6@*J?�    >�2�@�@�>m^�?8��?�    ?�w?��7?�H�?<8        ?�'Y>�� <�s`>�FI>��0?�?�?�X    @$��?��5    >�@�>am�>�ƴ?8�>q�                                                                                                L       parents[$l#L       =���                                               	   	   
   
                                                                                                           !   !   "   "   #   #   $   $L       right_children[$l#L       =         ����      
   ����                  ����             ��������   "   $   &   (   *   ,   .����   0   2����   4   6   8   :   <������������������������������������������������������������������������������������������������L       split_conditions[$d#L       =��u@?:0?ܭ��5^�	\Ϳ#�-�\��������V?�b@�Z����>�06�*�ɜ����>��D�����"*����<; о��_�9�?�DJ?�Ip�B�R>��P���о&[?l�?�C����(�X��>�"V?�w�V;���J��ꓼ�V
=���1���J$پ ����Z�<�9�ܸ6=�B���Y;�<�>�� @#�n[1>V���2�/ނ>�@��e�=��_�1�y>&ߩ=�.mL       split_indices[$l#L       =                                                                                                                                                                                                                         L       
split_type[$U#L       =                                                             L       sum_hessian[$d#L       =D=�=BzΕD-�TBF�6AP�|D��Bc'@d\A��BoU�D��@[�BUi�@��?��NB'��A��fD��A�<�?���?���AJ<B0Wn@[+@�p`A���A�x�Ay�7@QBjY>C�*?�ozA�U�@���@�ӎA
��B�3?��?�­@��?�@��KAi��A0��A2�@Z�AW�A��nBxC�~@� /@ ��A�C�@T/�?���@v�u?��M@��<@r%8A-��A�}lL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       61L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       5<]��=*҇�xhE={M8�h�W�0rʾ�%=�k����8���EW��cžֱ�>*k�<�� ;mu4��)��q��g�6��n�*}=H�߾��;��D�>P9�={�l�Ҥ��VJ�2[�=�.���;�>�謽ʭu=s����+�>��޾�Δ>ͮ�=��=�<־��=�f�8��>�\w��Vս��x?!Y�>V�辍K>��Q�ؾ�e@>��SL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       5                           L       idi/L       left_children[$l#L       5               	   ����         ����            ����         ����   !��������   #   %   '   )��������   +����   -   /   1   3������������������������������������������������������������������������L       loss_changes[$d#L       5@��@{|-?��@=�?�x?�@5    @#K8>���?��L    ?�I�?�?�f�?�J    >���?�L�?Y1J    ?�?h        ?���@5#�?�fo?ߔ�        >�C    ?#�?��?e��?�F                                                                        L       parents[$l#L       5���                                                     	   	                                                                                               !   !   "   "L       right_children[$l#L       5               
   ����         ����            ����          ����   "��������   $   &   (   *��������   ,����   .   0   2   4������������������������������������������������������������������������L       split_conditions[$d#L       5?+�>cV?��@$>���>IM|�=�A�3�a�QB�\ο]���Z��!&�-��:�y����ʿY߾o��+B<p�z<qپ�W�oͿ`�@�?Fu��g��V�Vs�#ɾZ���@�.$�9�Q=�q��Ĳ=���=�	<�ν�B���]��#�=�;½�5 ��_�>A�!=�¿���S==���{���<�=��1L       split_indices[$l#L       5                                                                                                                                                                                               L       
split_type[$U#L       5                                                     L       sum_hessian[$d#L       5DM#D9jB��D,��BF��B�RA���D)p�AI��B�NA.�GBMD�AJBCC�RC��?���A1��Al	A��@۾B1��?�p�A,X"A���C,98C��B�\A�"?�vC@l� A0�I@od#A���BQA.ζ@���A���BH�B�q�C�oA+��B�@@�-F@*>!?�y�?�Q�@
�1@�AN�A��A��A�?ݟWL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       53L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       c��D�>�=�C�2Eg��@O>*�̼b�ľ�P�<����<��|=��,>ͷ���֛>����ْ>�l:;��#>�P�6m���w�>V<���N��'_>v�$>��>�'�t3&<�e?"V=���<� b��7=����;������ؾ��H=r`��Z?�>�ad��6���>�g[>���?�ϼ��5>ӫѾ�WR���]>��ټzO�>�S9?Bp�>-?S��L]�^��>��;n��>�u��z.�>.�`�>�v0�N����>D�!�Ѿ�P�>��V?8�(=�z��KxH?!�y��=��>�{B�>��E>�X=��=>�>��K>�LC�M�l�����8VU�xb�>c�L=Ӄ? ���>16�<c��>��N?[�>s`�>��.�FpL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       c                                                  L       idi0L       left_children[$l#L       c               	                                 ����   !����   #   %   '����   )   +   -   /   1   3   5   7   9����   ;   =   ?����   A   C   E   G   I   K   M   O   Q����   S����   U   W   Y   [   ]   _   a����������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       c@��1@�b@F@ڸ?� �@1b�@�?_��?i��?P�P?6�?�e�? �?�C:?�$q?`��    ?\��    ?8@�?6 ?V1�    ?���?�`=�Q >���?�;�?`M�=�� ?[?��    ?]��?_�?/ �    >��`<��>�>r"@��@��>�q?��>ָ�    >���    >q�0?��9?�o?��]=�H�=a�?7f                                                                                                                                                                            L       parents[$l#L       c���                                                           	   	   
   
                                                                                                               !   !   "   "   #   #   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   /   /   1   1   2   2   3   3   4   4   5   5   6   6   7   7L       right_children[$l#L       c               
                                  ����   "����   $   &   (����   *   ,   .   0   2   4   6   8   :����   <   >   @����   B   D   F   H   J   L   N   P   R����   T����   V   X   Z   \   ^   `   b����������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       c��(�5 ���о�q@ n��:2�@��@-믾�p��+�����>~|<��>]R@,$���=��F���>
��w�z@�}?�!���5������vih�%[�?��>�sR��F?
X>9g�>Y~R�u�>�U�?�:[@y��	D��/,@N{@�3�Z@��g� �ZR>�8��!Uj���z>#.,����=�b?�@^<��h;�K?�;�l�>��Y@Y�'��[����=�=�:�`�=�Yܽ�=(7U�3@�>���x\S��Q=���B=b��a=�u�>]y�<��t)�>A����g�<�K����=��>�<��<d�>~�=����v��M��]4g��=��.<.��>��*Z=T��;��=�A�>�gh=��=�J8�n L       split_indices[$l#L       c                                                                                                                                                                                                                                                                                                                                                                  L       
split_type[$U#L       c                                                                                                   L       sum_hessian[$d#L       cC�Z�C:�C��(B�S�B���C2TC��A��B��YB�)<A$�B�!B�AB�A&A��PA��J?�y�B�J@xA�AW��Bhn@�ŭ@#%B���B#&#A��A/ B�B��@ρ�A/U�@�.A�BO$�A��A	�@���B_}j@
�@<��@,��A6nBS��@�ZBz�A#�A�e-@��@D��A��]A���A"ٰB}!�@,;o@r�EA
�?�Y_@+=V?��B�JAT�%A�\A/�@١�?�^E?ؼ�BX��?�L?�K?��9?�Q?�X�?�ĳ@�O�@û9A���A��%@�H�?�E�A��AX�p@x�H@�٪?�;@���Aa9�@���AI

@�C@���@�fB�oA��?�:�?�<7@*�N?���@�8�@��L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       99L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       7;�u?�׬�=�����-�<�3�>����;p��� ����o��ݫ<�h?>��>�V(>�u�;�k�b���R��Mi=��p>GR� ��K*�>�?=Ś���>n���o���<��=c"'>�z\�R�W>�=�>�J&>�Ց�<g���E? �2�4h� ѹ��69>yǰ=��K�D��>�t�=���;��)��	�M>���>�kT���L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       7                            L       idi1L       left_children[$l#L       7               	      ������������               ����   ����            !��������   #����   %   '����   )   +   -   /   1   3   5����������������������������������������������������������������������������L       loss_changes[$d#L       7A'u?X=�@#��<�T >���?��5?^�l            ?�?�#&?�?��>�LX    >CW�    ?�g%@$"�?�sL?d�        :�(     >�-�?�B    ?�.�@��?�Xi?��(>�D�?��>�!I                                                                            L       parents[$l#L       7���                                               
   
                                                                                                     !   !   "   "   #   #L       right_children[$l#L       7               
      ������������               ����   ����             "��������   $����   &   (����   *   ,   .   0   2   4   6����������������������������������������������������������������������������L       split_conditions[$d#L       7��u@?:0?ܭ�@A�����M蔾��_�  �󚿾�2?p����6�� ��4=���?@1¾� ?���#cx?�	>�06��4�s�/�3�L<�̾��V?���	�v� M�?�z?U�/?��>�"V�Q��?���>�a� $1;�0��!�>L���}��E���=��7<�C��l�>��=��;^p�e�%A*=�h>s��(��L       split_indices[$l#L       7                                                                                                                                                                                                     L       
split_type[$U#L       7                                                       L       sum_hessian[$d#L       7D5�BQ�D'�/B!�	A@ևD�BN&�B��?���@0��A��A��D
�ByA�2l?�@�@���A�aA#1C�iEC���A�6?�+�?��>A�X?�Wr@�@�M@]��B YCiJsC�X�B�q@�~�A�h�@�5yAK��@g�0@7t�@��#@+�AӦxAQ4uCH�B�CC�R�A�]JAd�hA��/@>�?���@:W�A��@7l�?���L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       55L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       9<Rd�=6���>=?�����I�3��?�=`ｾ�����U��xJ�l�>��w=�-����߻C����4�>B'�2Y-��i]��|j��s�����?rw���>�:b�=��Ӿ�����|���D�A�>��Ͼ�G�<�U���ǾF�w?
���Gپ���=-0�P�>I��>X,�����|�?��=/��j����>;|7>��о�F�����k>#�6����L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       9                             L       idi2L       left_children[$l#L       9               	   ����                        ����         !   #   %   '������������   )   +   -   /��������������������   1����   3��������   5   7����������������������������������������������������������������L       loss_changes[$d#L       9@���@J��?A�0@ ��?&�?k    @o2>s�>���>���?xG�?>`@@$�?���    >L�P>�>Q��>�~8?�r�?;n�            @Yp�?�u�?���?t�                     =Ʈ�    ?�        >�O�?H�$                                                                L       parents[$l#L       9���                                                     	   	   
   
                                                                                       "   "   $   $   '   '   (   (L       right_children[$l#L       9               
   ����                        ����          "   $   &   (������������   *   ,   .   0��������������������   2����   4��������   6   8����������������������������������������������������������������L       split_conditions[$d#L       9?p]�?8�?��@$��?�*F���?΄�3�a?��|>��>����Sˠ�����#v��j�s���ʾլ��f�?��f>�X�֡���&>(�\�����7־�n�& ����6���#�"=��,�߉(?b]l��޾��K>%��^O?���?��>�y��=rS(=����0B�䕊>3��<7��ӳ�m�=`�v=��`���4�v��t=D�A��C�L       split_indices[$l#L       9                                                                                                                                                                                                                  L       
split_type[$U#L       9                                                         L       sum_hessian[$d#L       9DD�eD8��B=֮D0�ZB�Bc�A]̵D-�A@�@@�{8A�U)A� @>/D�PB���?��jA)��@[t.@��!A�� @ń#A��A"�B?��?�Q�C��C�K�A�K�BU_A��?�).?��-@+?�Ȣ@��ANoU@���?�[@�L@�AN�%B��Cn��Bx�Cn9�A��j@d\bA��A�,X?�1�?�
?���@�N#@(1�@�~�A%؀@$�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       57L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       ]�˼��/�S=���%侹�=�$�ï!��}<�7�в�<w��=c�>h.�'5>�-Q��J >&>��ݼbFj�-�����? �����P>���:�L�>��3>����lM��	=?�ҽ��Z��8�헒?%'�{7��R�<�:�=ë������8�=H�����d=�Y�UX&?!������=A�,>8_�����<xdG���о���>:�;=�P?�	�T��=Ƒ�?IΏ=��O>+|X���O��8�=�
��N�>���=�� �=鼿 R{�6�"=�Y�>O(�����u�>�$?=0J=E>!���� �=�����ݣ=�x>��<.#��tʾ��Z>��L�ņ��D�=�}���>����!�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       ]                                               L       idi3L       left_children[$l#L       ]               	                                 ����   !   #   %   '����   )   +   -����   /   1   3   5����   7����   9����   ;   =   ?   A   C   E����   G   I   K   M   O   Q   S   U   W   Y   [����������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       ]@Ī@�C�?�4c?�,?�K�?�>,?��!?0�?p�d?>��?%�?�	�?���?��S?��>w=     ?ͽ3?N�X?3t?%�p    >�t�?�5?��(    ?���?A,?���=��P    =�T�    >��p    ?7�?E[�?i*?7l>�H@<Ԇ#    >�1?i�>�zh?u�?r�|?�s�>*��?>�h>�-�?\��?<�                                                                                                                                                                L       parents[$l#L       ]���                                                           	   	   
   
                                                                                                         !   !   #   #   $   $   %   %   &   &   '   '   (   (   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4L       right_children[$l#L       ]               
                                  ����   "   $   &   (����   *   ,   .����   0   2   4   6����   8����   :����   <   >   @   B   D   F����   H   J   L   N   P   R   T   V   X   Z   \����������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       ]��(�5 >!j�4 @ n��sb@��@c���^p�+��@Ij��p"� i>��#?�0���=7�a�4�޿H�Ծj׳@�}>S,���^�fyT�l��>��?���=�{�?6^��༮���^���%�!sݽ��ܿT�>4'Ӿ�'?��T�/,�cQʽ��>�Ӭ�o<���<lgA���G?���>���T�@
���c`@�=�0>3ǥ�6�<�H�>r+=�c=M�j���,��w=>��+_=íھ ��=P4�c�I����[9�=i=x�1�����&�=6�>c�<l���#'�A&=!0��=+=H>&S;P���&���m=�+�����R�=�K��=�����[�L       split_indices[$l#L       ]                                                                                                                                                                                                                                                                                                                                               L       
split_type[$U#L       ]                                                                                             L       sum_hessian[$d#L       ]C֫`C*S�C��rB�E�B�a�CN:HBS"nAkTPB��RBw��@�AcB�MB��DB9� @ˊiAUպ?���@��B��AF�QBFG�?�x@�c^A_�TB՚A���B���A�{�A��@�?��J@ �A1M�@��@QCA!��B�W8@���@���B=��@��@�8@���@�ZV@��RAv��B�ɮBuN�@��@�i�A��%A,IyAk��?��d@W��?�<�?�N@M�?��@�@�ϐA���Bd@�@S_�@�C�?��H?�rB6�N?�xC?�|@O��?��1@A�@�͒@���?��@Ȝ�A4=Bo�A�'�BA��AND<?�iN@Q��@ ��@4OPALk@Ux@N�9@�LVAQ��?�sL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       93L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       7;w���c�=�ʾ���%���]�=��̾��\�fվm�=��R��b;��3=`��>�GZ��.�=�����$_>�[a=K�0�4 ��0~�=�������������>��;�3L>�0`������>����Q%>殯=����ݭQ��>�s;�de����<═�~�>
�=���>�O�o� >[�0�_��??>=
�����h�?0� �B=�j*L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       7                            L       idi4L       left_children[$l#L       7               	      ��������   ����         ����   ����   ����            !   #   %   '����   )   +   -����   /   1   3   5��������������������������������������������������������������������������������L       loss_changes[$d#L       7Am.?@�8@L;� >�)�@k�@&O�        >/��    ?ڮl?���?�D�    >#i�    ?Q�    ?���?�b�?�4?�v:�B >�0�?<x(    ?��F?��?��    ?S�?�?��@��                                                                                L       parents[$l#L       7���                                               	   	                                                                                                           !   !   "   "L       right_children[$l#L       7               
      ��������   ����         ����   ����   ����             "   $   &   (����   *   ,   .����   0   2   4   6��������������������������������������������������������������������������������L       split_conditions[$d#L       7����?:0>�]9@9R?v��U�*@���%��*��@ ��=W2@=�D>*X�H�'>*�>k�-<�t@'�>�n?)�@Z`�l���@>̾�&�?nm
?�C6=΋O=3k��Ž�>�.�=t9�x�ĸF=�PH�0c����m=�Wý�EF�袥<�W�"�`=%��<�Y>�c���=�ꄼ�K�>2�=����V˼���>T#4�h�<�fL       split_indices[$l#L       7                                                                                                                                                                                                     L       
split_type[$U#L       7                                                       L       sum_hessian[$d#L       7D."�B.�zD#5�B��A-wCBȃC��A�	?���AQw?��B/�?C�sC��A_<�@�CN?�~�B%@)�oB�A��B�5C�pp@�BT@X�B i<?�ہB�QA�	�AϮ�@i�@���A�kA%T@C�E�@K�T?��?��@fB��@��BK^BT��AtaA��A�ד@�]u@+��@
@�rnA���@d@ؤrA�/jC���L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       55L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       C<._�=>{5�[�=vTK���޺ؼ��q��=��Y���D�?~��U��q�={JĿ"�N�H�+=t�>�K��ӕ=��1�⡿=]æ�{����K���i���=�a�׉%>剼�c�?>#� =,w?���Im=�����|>�=��Ϳd����>�R�P
=�=m?�s� QS�����ߪ>]x��a�=ߎ?'�=��i���˿]�<.g1?�>�����.�<Wȿ$+�>�b�?���8}<��ݾ��ĞԾ�/�>K�$L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       C                                  L       idi5L       left_children[$l#L       C               	                        ����            !��������   #������������   %   '����   )   +   -   /   1��������   3   5   7   9����   ;   =��������   ?   A����������������������������������������������������������������������������������������L       loss_changes[$d#L       C@��C@(�v?�=?�?��?�(�?�?�?�4�>�x?r��>8�>7}8?��3    ?�~x?�i�?�H�>֝x        ?d��            =�?�v�    =�/P?t�|?⌄?ĳj>���        =�+@>��?Y)<	t     ?�V ?I�        ?�A ?'�                                                                                        L       parents[$l#L       C���                                                           	   	   
   
                                                                                       "   "   #   #   $   $   %   %   '   '   (   (   +   +   ,   ,L       right_children[$l#L       C               
                        ����             "��������   $������������   &   (����   *   ,   .   0   2��������   4   6   8   :����   <   >��������   @   B����������������������������������������������������������������������������������������L       split_conditions[$d#L       C>:	?g(>BY"@j�Q#t>�n>2�=�&W=� 5D?��2�!�X?���C�>�%:�#�-> xV���<�Wվ����������k��8�����g֨�RJ���?�$��!&�!sG>(�н��<�g%�<����"ξ��ǽC�?@1¿�C�=�>4����@�+���3=���2+<=r�>I+Y<�V��'�pJ;QH�>9��=�N����b�E:>+�e���<D���ռ��̾O�=tĒL       split_indices[$l#L       C                                                                                                                                                                                                                                                   L       
split_type[$U#L       C                                                                   L       sum_hessian[$d#L       CD=9`D��C�IDoTA�5Bv��B���D��A/ezAm�	A�b@�ӔBZ5^@ʪ�B�	�D��AG��A�+?�b{@���A��?�1�A�0?�@��PBH�+@�)�@�B�4DB�}Cކ�A+�?�p&?���A��@6��@��@��K?�$A�K�A�Tv?�Oz?��Bj��A��A���B�^O@C�C���At�?��3?��@��?��]?�ב?��"@��?��%@EA`P�@��+@W%A�o�@�BK��A��L?���L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       67L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       [���+���L=�o���;���>�1=Y��<|���0����3<�=���<7>��<��>� N�6I>�yO��]�=yz��!��-���&>�p��s}j>j�TS>�ͣ�)կ=�1T?Oy�>)�=g���N�=[��>��E���!E�>���aŒ:3^"���d���u>�>:>`�\��W�?D�T�� ɾ��=�C�>��~��Ju>�a)�"�ٽĺ@��
�>Iq$�m�>Û����Z;uN�>�Go��m>G��>�3��$�=����%���L>�� /P� �S>�m���2B>��[��N�k���-=d->��6>�I���f�R	�>E��?=�=�}>�����>�l� ���7�Ź"L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       [                                              L       idi6L       left_children[$l#L       [               	                                    !   #   %   '   )   +   -   /   1����   3   5   7����   9   ;   =������������   ?����   A   C   E����   G������������   I   K����   M   O��������   Q����   S   U   W   Y��������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       [@��@�^?�S�?�R�?�Pp@)[?��?�@u?�]�?N�`?��=? �>��`?��?�q{?t��=�N >}Z�?���?!��?=�`?�z?��g>_�j?k�    >�P?~$?���    ?�?�5�?��            >�}     >��?��=ma     >%�            ?�>��    >h��?3�1        ?a�    ?lL<?@�b>�Ǟ<}[@                                                                                                                                L       parents[$l#L       [���                                                           	   	   
   
                                                                                                                             $   $   &   &   '   '   (   (   *   *   .   .   /   /   1   1   2   2   5   5   7   7   8   8   9   9   :   :L       right_children[$l#L       [               
                                     "   $   &   (   *   ,   .   0   2����   4   6   8����   :   <   >������������   @����   B   D   F����   H������������   J   L����   N   P��������   R����   T   V   X   Z��������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       [�%Ʉ<�h���B�>G��@ �?��@�?'~�?s��@�?��>��6����?\Kb@��6����?�~�?��k�/�=Х���@���ë�Z�N�(e1?�ڌ>��;>+��>x�{?�j�?N�^?���<���>��� Gz�3�r>U׿�����6>z���Z���=�ƞ��>kՙ?5�J�=^�<لO�m�;�>�C
���1��9��ν�>^�>�Ӭ?�	:�/0>�v�5�=o��=5,>��Ņ<���������K�=���`�m1>���o�=�|��ϑ�������<���>�=�$���Y��|�=mWq>�=��=�6t�*W�>ۼ���^C��D�L       split_indices[$l#L       [                                                                                                                                                                                                                                                                                                                                        L       
split_type[$U#L       [                                                                                           L       sum_hessian[$d#L       [Cʝ�C~�CXJC>̥B�-�B7H�B�%C((JA�"�BT�A1b[A��A��B�<�A.{C"@Å�Ak @�O&B@U=@�m`@��>@�y@�7�A�?�LA�1�A�x�B|�9@Dߞ@��dB�*�B��?���@�Y�A2��@a�t@$�;@�։@-wPB5}�@�,@)J�?�p�@�@d�@W�<@���?��,@��2@�2�A�A?��3Aͺ�@��Bq�A̖�@�X�@
[�B�x�A%��Bm xA�P?�F�@�+@�@@?��t?��,?��B0�*?���?��F?�!�@�y@<|"@,��@'�u@B�?�Bs@4��A�z@ڕZ@�]�A��u@�TfA���@��o?��?�	F?��
L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       91L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       5;�v����<�+"��Lw��T<R�>e6��^Ŋ=�|���<�������>�Kv����;oZ����4>~�v�ak<��>̛۾4)�>9u>������
��
�>n��x�Ѿ󝪾�7=�W�?M��<�w=`��n=Ë�>��A>+y�����~5>�IL�N�<�DB��w(�؈y>�q徱�R����=�y~�2�>�n����>��gL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       5                           L       idi7L       left_children[$l#L       5         ����      	      ����                     ����      ����   !   #��������   %��������   '   )   +   -����   /   1����   3��������������������������������������������������������������������L       loss_changes[$d#L       5@ӫ�?6��?�R�    >V� ?�)�?M >-$    ?> 6?� ;?v�U?*��>��>z�E>��    ?)�?�U�    ?J�->�3�        >���        ?s{�>�
h>֘h?��    ?���?,s�    ? ��                                                                    L       parents[$l#L       5���                                               	   	   
   
                                                                                               !   !   #   #L       right_children[$l#L       5         ����      
      ����                     ����       ����   "   $��������   &��������   (   *   ,   .����   0   2����   4��������������������������������������������������������������������L       split_conditions[$d#L       5����?:0?ܭ���{?v��g�i�T�z?\�8<��Q?�g��Yf$�h88;�A:>����i>��B�r=��z?b�X �=���>�9�?��P>w���=�u{=�Y'��3�?T����V�6�?�$z>v��?0\�\�{�*�z����>_[=M6+�Ĵ��d@=ξ\�(^d<(��
���|>w���0c��)q<��˽V˹>u7��d�=�>�L       split_indices[$l#L       5                                                                                                                                                                                                L       
split_type[$U#L       5                                                     L       sum_hessian[$d#L       5D(��B�D4jA���A"p�D��B8L�AV?���A~x�D��A<�^B	�@��:@��Ac��?�y�A��D
u�@K%�A	��A�cdAE�I@Cy�@4,�?���?��@�:�@��Ax9�@���?�p�D
!@�O@�GA��<@�Ġ?���?�_(@���?�@���?���A�-@��[@=�@!��C��.C�@�G�?�O
A!�@�,L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       53L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       C<��<̱?��x�=�@�}��=O����.�=I�8�1�K��r��A}>�
���nϾ��7>9�>~z=�ɾ��f�Ļ���뾽���Q�8>����NV���G��_���1&> ��>��	��T3=(�'�B���>$ag��֪���.��̼=�/���k>�;�;z�k�Ȝ.>�e�H�Ǿ�N�>p\��9�=���?��!,��)&�=F���wu5>��ǆ+�M-�D5��g>Թ�����>:���.?'��=�����m��
.��.L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       C                                  L       idi8L       left_children[$l#L       C               	               ����         ����            !   #   %����   '��������   )   +   -   /   1   3   5   7   9   ;��������   =��������������������   ?   A����������������������������������������������������������������������������������������L       loss_changes[$d#L       C@K^�@�9?��L?۞*? <?Ow�>�)�?�Q#?��<?��    >/�;Q� >�Ȑ    ?���?���>�xX?���=~5�?h�    >*Y|        ?Z�>�(�?���>�N�>�K�?���?1{=�� ?Ý�>�}�        ?Z��                    ?�w<��                                                                                         L       parents[$l#L       C���                                                           	   	                                                                                                                 !   !   "   "   %   %   +   +   ,   ,L       right_children[$l#L       C               
               ����         ����             "   $   &����   (��������   *   ,   .   0   2   4   6   8   :   <��������   >��������������������   @   B����������������������������������������������������������������������������������������L       split_conditions[$d#L       C?�2?g(��@�> ݼ@/�@l��j��@,-��QB�����п0�8���=_�m��i�{��"�?�{��e�n>���{��>�Ӭ��ν�#>�"��@�n�h�|��?7��?6!v@<>��P��'@S���Ȟ��>>�<��>�@:�t���k=��>�N?��M=�k���<�*�>2:W�Ah��J��<n<s��y�=�n��mξ�нks񽙊>=�E ��Y�=`Y'�P�A>I:e<��s�C���,t8L       split_indices[$l#L       C                                                                                                                                                                                                                                                 L       
split_type[$U#L       C                                                                   L       sum_hessian[$d#L       CD7��D.DB�D&�!A��_@�@�A�~�D�B��A�gA��@��C@�pA��f?�g�B'DcbAj%�A�@�3�Ae�	?���@��?�L/?�r�@���A�3A�PpAG�0@��Dݮ@I�A7��AI�rA`�?�ɋ@��&A;݄@(F@E�?�� @=[L@�J@A�bpA��@�٥@Az:A��@�T@��DN�Ac��?�<�?��A	�@;x@@���@��@�	?��A*�x?�]@Cx@A�A��?�&@L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       67L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       G�� ���=����B�᾵�;��l>۾�l:ny��ې<gڻ=LGq�J�->���=��.��V�=��y=����@���ر>*�v�b�\>i�<�}>�ᾪ�[=5�l>w=���������;�?w>���t:=T��='p�>bk����>��k�U��=(���	�T?�-=�(=�X���Ѿ�b>9�E=bb�>�I��o��>]\�>�o張R3�� ���W���R������+l=İ&>*)?1���=.>�n����C>g�C�֗W>�I���OL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       G                                    L       idi9L       left_children[$l#L       G               	                        ����      ����      !   #����   %   '   )   +   -   /   1����   3����   5����   7����   9��������������������   ;����   =��������   ?����   A   C   E��������������������������������������������������������������������������������L       loss_changes[$d#L       G@��k@M�"?��3?�u�?�N�?�3?�?0>��?���?��??c�?KY@    ?��.>�~�    ?��h>r��>�z�    >���?��?G�>F��>�J�?��?���    >i�    ?e+�    >S��    >xW�                    ?=BZ    =��         >���    >���?K�\?���                                                                                L       parents[$l#L       G���                                                           	   	   
   
                                                                                                   !   !   #   #   )   )   +   +   .   .   0   0   1   1   2   2L       right_children[$l#L       G               
                        ����      ����       "   $����   &   (   *   ,   .   0   2����   4����   6����   8����   :��������������������   <����   >��������   @����   B   D   F��������������������������������������������������������������������������������L       split_conditions[$d#L       G�Ke�<�h��1����@5
��(z���@c�?U4@XT����@�?Ky�>��?���<���?��@@;&�=M2�@�>X=ҾZ��@7쿅>�?O��?��ھ�o���}�����^p>��?�þ<�{@2�<H��=��$���j>H��S˿:Z�%�e?O��=��<�jK@���B}=�6�>� �@D����(=��@=�쭻ٕ׾f��ٛ��u2���+��4<��=L �>U����~<48>(��h�=��)� �5>	ƽ���L       split_indices[$l#L       G                                                                                                                                                                                                                                                            L       
split_type[$U#L       G                                                                       L       sum_hessian[$d#L       GC���C y5C_�B�TB@f-CB��;AoͯB�şB��A�eBܒJA�W�AJϰB��EAZ�i?�Z1B�7�Ap,B{K?�)@w�[@�`B��0@�Q�AfM�Aa�B��@pja@ 6�A2t�B�>@�ո@�C?�pSB�P?�?^?��2@5p�@=�g?��B�A�?���@/��@�v?��AU˻?�}�@ң�B^�"A�W�?���?���@�f8B�C�@��r@��B��?�3HA��B��p?�+�?�-�A@J�?�	�@$�@��rA�V�BP�A�jG?���L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       71L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       1;y]ھ�x�<�;������<.�>U�����L��⓾��<�M%>�
>���>�l��'O���3��|<eu>�꥾$>RSu�r��>H�8>Bvξ���xX�<��+=��d>��>hċ��5ϾA�X>Ꜿ�ˏ�1!z��>�N����E>��?Y�<��l>�k+���E��V��c��y<=���>"�v>�LL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       1                         L       idi:L       left_children[$l#L       1         ����      	   ����            ��������   ����                  !����   #����   %   '��������   )   +   -   /����������������������������������������������������������������L       loss_changes[$d#L       1@�U7?:JH?�V8    >6�j?�?2U�    >��G?�;�?���?-u�        >��    ?p۴?���<�.@?K�?�>+�    >�t    ?.��?���        >A�+=�X>G�>�V$                                                                L       parents[$l#L       1���                                               	   	   
   
                                                                                            L       right_children[$l#L       1         ����      
   ����            ��������   ����                   "����   $����   &   (��������   *   ,   .   0����������������������������������������������������������������L       split_conditions[$d#L       1��u@��?ܭ��<�����M蔿)B>������2?p��@7��?��>ڨ=��j?v���?���gvԾo��>�q�\���=p��?��� HV?�g��aF4=0p>
p�>�.L@$�H@/�=�9����T���'�e>������=���>,;��O=����� �sμ�u��^I<��f=CP�=�(L       split_indices[$l#L       1                                                                                                                                                                             L       
split_type[$U#L       1                                                 L       sum_hessian[$d#L       1D#�sB�De�A��FA.ŽD��B,p�?�d�A�&A�,�DU�B$i@�a?�"�@���@�V�A-�D
Ʀ@�n�@�*wA�>5@�v?�,v@��T@6�A]��DO�?��@��B@(�M@_��@-�AٛZ@a �@G;�@s��@.4AJ�,?�C�@~�jDQ&?�	?�W�@o?�k>?��?�:A��A/�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       49L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       ;;��U=���q=7 ���QR;@�h�SZ�=Qد��B`=臢��oϾ�z�=�ſT�*e9=3<>�����!=�~�چf�������vC=����>��=�E�k<�$�>E��>�q׾�=��
��y�����1�<�)>�ç���J���\?M�뾖�����p��M�=I�'��>���YJ>�n�?7竽�����=�	���9??�W���O�=��(�$q#���&L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       ;                              L       idi;L       left_children[$l#L       ;               	            ����         ����            ����������������   !   #   %   '   )   +   -   /��������   1��������   3   5����������������   7   9����������������������������������������������������������������L       loss_changes[$d#L       ;@%��?�H?��?�]v>�z?��?���?��>�ۀ    >�>Ap ?���    ?��x?�\?���>��\                =�' ?��T=Z�@?��?S��?���?�f>�^�        =�D         ?�%=?�SY                ?�?T�p                                                                L       parents[$l#L       ;���                                                           
   
                                                                                               #   #   $   $   )   )   *   *L       right_children[$l#L       ;               
            ����         ����             ����������������   "   $   &   (   *   ,   .   0��������   2��������   4   6����������������   8   :����������������������������������������������������������������L       split_conditions[$d#L       ;>:	?��|>BY"@j�Yq`>�n>2�=�&W=��a=���
�!�X?�n\�6�Q>�%:=X�4> xV���<����q���M��8!����ͨF=�+�� g>��� �>�x�m��J
<�Js�<��)�̼���T��>AA��`� O8>vܴ��̞�Ұݾ��T<qE#�Io=�7���_�=�T>\������;t<�>۾"Y>;X|��[5��_�<ʰ1�ET���L       split_indices[$l#L       ;                                                                                                                                                                                                                      L       
split_type[$U#L       ;                                                           L       sum_hessian[$d#L       ;D2��D@�C=@DC�A?+�Bf�eB���D�#A��?���A+�@�K�BL��@��cB�MD�KA<��A4$?���A�?��?�:@���B;�U@�L�@ �pB�FSC�TMB+�LA"�^?Ь?���@�G�@yq?�	�BIA-�2@@�O?�;�?�u�?�7B"�A��gC��B,!�BC}@��w@��@��-?��@��lB@.��A ��@3�qAW��A�{�A�ziAN��L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       59L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       C��n(���=n������m"*=� �����=�"��Q?=�m�(�E<��->"S����=�W@�M�d>����۳<5�-?�1=KĘ��h��w>r���>H|C>��)=�k2>��꾉j�><����@���%?��b��u=�꾾��>���K>_�	= }G�t>>��=����>%:��b�>"i���>�r";o$��Է�c��?\��2A�>O��;����x>�0<Q>�'�>�x���IL> 3@>�Ӵ����>�cj>"c&���L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       C                                  L       idi<L       left_children[$l#L       C               	                        ����      ����   ��������   !   #   %   '   )����   +������������������������   -   /   1   3   5   7   9   ;   =   ?   A��������������������������������������������������������������������������������������������L       loss_changes[$d#L       C@J�d@/t'?|Is?vEh?���?~��?$\�>��>�= ?��?b,j?�2�?���    >�^>�`�    >K��        ?E� ?���?M�?�K�?�    ?v2�                        ?-sz?^5�>�Wh?N?��>�%9?Qd�?��>�l�?{�@?f�                                                                                            L       parents[$l#L       C���                                                           	   	   
   
                                                                     !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +L       right_children[$l#L       C               
                        ����      ����    ��������   "   $   &   (   *����   ,������������������������   .   0   2   4   6   8   :   <   >   @   B��������������������������������������������������������������������������������������������L       split_conditions[$d#L       C�Ke���q??�ȿQ��d��1��?��=�Zx@���w�#?1��?&)���ѾeD?�tN�6�=��?�y;Z(7>-�;�J��@#��@����'>���>�?��=�����=b>��
�P�Y�:�ܿU����?�|@3���䉽ۋ?��|����?y��?���@D��;'=:)K��[=�U�:,���ռ��&>.o4�U�=�:�aI�����=��;z�o>�>HU���=@=�>�l��E=��=B�a����L       split_indices[$l#L       C                                                                                                                                                                                                                                            L       
split_type[$U#L       C                                                                   L       sum_hessian[$d#L       CC�>CUdCX�B��B�JCPe�A6r@�ۿA�sBW�B���B�v�B�T�@��O@CY*@.0?�d�Aռ�?�a�?�m�BRǤAߐTBVBͼ�A���A)-B�/?��D?��?��@?�z A�"�?��@@�tpB9�A���@5��A�2@���B�}�A��pA���@��B�hQ@��@�@��mAc��B �A���@y"�?�g?�m@�w�A�zE?�&	@p �B�s�@���?�+	A���A0�~@��@WO�@�c�B~:Z@��;L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       67L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       A;��;���<�:��ʥ�RL��E#=%w����W����x�t=��J=�y>��>��T������ʾ �+>�p��v=;u������:>��Z�q�1<ݏ��ž<K���">�E>؛����=������<���>+O��� =m�(�ͭ�>��>�n=<,���7<�AM> s.��el�_���<�3>�>N�}D ?	�>�Q����~��V�>�t��cw=���o�4<�e>y�E������֨��B��>�_L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       A                                 L       idi=L       left_children[$l#L       A         ����      	   ����               ����                  !   #   %   '   )   +��������   -   /   1   3   5   7   9   ;   =   ?����������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       A@��'?-0?�o    >p�@(��?���    >�l�?��?��	?��?BCd    >�=x9�?�(�?�g@?pi?׆�@�?"�4>+_�>m��=���        ?���?} ?� �?���?g4�>�h�?��R?��?N0h?�*                                                                                                                L       parents[$l#L       A���                                               	   	   
   
                                                                                                                       !   !   "   "   #   #   $   $L       right_children[$l#L       A         ����      
   ����               ����                   "   $   &   (   *   ,��������   .   0   2   4   6   8   :   <   >   @����������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       A��u@���,�������?^�9@���֙���2�G�?�3"?�^=�7N=�:̾��V>�zK>�%>�JA��?^�&�:>��R@%I?G��>�8��?��a�>� G?!gϿf{�?�*��"*�=��ֿQx>��?*�4?�߶���_=�AM>�v<H5��v;�*=@�8�p�>߼1�;�Wq>%b����>�_=�.�� W���=�%����<������<�4=���0��6|ʽ ˃�i�j=.�?L       split_indices[$l#L       A                                                                                                                                                                                                                                      L       
split_type[$U#L       A                                                                 L       sum_hessian[$d#L       AD�_A��-D�A�"pA%�yB�1�D��?�)�A�?B=ѿB��C��,Agsx?�0�@�@SAjIBP�A���An�C�+B�!@JܒA4�S@��=@�-AG�@D�A�AlA8��A���@�[A��@�ȐC� B���Ap� A���?ߓx?�%�A#L�?�|�@/Y�@T�?�)[?�z�A�A4��AA@�h?�Aj�@$V�@�x�@
RM@Ҷ~@�&f?���A���C�$B��A�|%A*@�˫?��HA���L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       65L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       ?;�Y�<��z�k<�M��W=�J����c=L��"�ѽ��@���>����k���yA>??�=����D�������˳���<�}�S�ɾ�>B>%��<�^˾ܱ�;��<����>F������C=���>"������s-=����A=��ߖ>�_=����%�>B�1�=���?P���()(>�Tz��Tw�N�K��i�{>�n�>T6P������/��熀<�|�?-�K<��ݾ��>�-��m�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       ?                                L       idi>L       left_children[$l#L       ?               	               ������������   ����                  !   #   %   '   )   +   -   /   1   3   5   7����   9����   ;   =��������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       ?@{??��k?Q-�?�kc? N>�S0>��X?�l�?i��? ��            >��    ?���?�gR>�l?_��>��0?-%?f�}=��@?���?^?q�r?�|z?��>� ?���>�"v=h-@    ?0�;    >�l�?.Z,                                                                                                        L       parents[$l#L       ?���                                                           	   	                                                                                                               !   !   #   #   $   $L       right_children[$l#L       ?               
               ������������   ����                   "   $   &   (   *   ,   .   0   2   4   6   8����   :����   <   >��������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       ??�2?g(�h�@�> ݼ?�@^@y~@,-���N��=�[��L�>$�=e�=6Z��3���"�?�{�?�>���"Nv?�T��r>�z�9��-�@<@!�'��'�(2��YM�<��>�����<��>$v �����=�2<<cl��i=h�9�UE�<��>z�Z�I��=�����2)�U+�tx���IJ=��=~����)���׾
�M;���>P��;���:�=�6���EL       split_indices[$l#L       ?                                                                                                                                                                                                                                   L       
split_type[$U#L       ?                                                               L       sum_hessian[$d#L       ?D/3�D&�B'=D �A�~�@���A�b�Dt�B�:A�M�@�Á@P��?��A���?�A�C�VC��uAUx�A�N0@�~�A.�jA^=�A[��B�U�C#�2@�('C���@2�A(��AAL�@���@��?�s`A	�@��A�L@�1?���A@��B�OrBl�B�-B#��@X:<@?��C�%I?���?�|@�E�@yC\@�O#@�I�?��[@ս�?�
�@��s@� ?�c?��m@��@1��@�mL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       63L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       Y���S���=��ͼD����$>6�]��T�<��*�Ri��u+���q����>}뾬D�=%��1 �>�=����=2⹽�#3��[�;P���ޕ�@�z=�=	>��=����=��>�wj<
=H趽��,>�2����=���ȼ�'%�>�uྃd�>ۢվ �U>~4���yK>Eq�>�>��4V=���>��=:�?��=�P?�[����=��Z<�B?]��1�>\_�?Hb���>Q�־��v>���4���dK=��>@o������t�>cl��	�>�>�cھG!�����>�2=C�6>ཪ>��_��R�>��R�A꫽}N�>�Qc�����Q?0��<oUgL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       Y                                             L       idi?L       left_children[$l#L       Y               	                                    !   #   %   '����   )����   +   -   /   1��������   3   5   7   9   ;   =   ?   A   C����   E����   G   I   K����   M   O   Q����   S������������   U   W����������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       Y@,�6@OK?��?��F?��?{�?l�?�_"?#�?X�@?;��>�:?}�0>һ�?1}?2+�?�R?GH?@�\?Wn�    ?Z�    >��#>��>��?S��        ><4�?�|?��?x��>�{�>���>���>�1�>�0�    >�=�    ?{9�?�$p>ә�    >`
x?@�>���    ?W^M            ?}d?�+                                                                                                                                        L       parents[$l#L       Y���                                                           	   	   
   
                                                                                                                 !   !   "   "   #   #   $   $   %   %   '   '   )   )   *   *   +   +   -   -   .   .   /   /   1   1   5   5   6   6L       right_children[$l#L       Y               
                                     "   $   &   (����   *����   ,   .   0   2��������   4   6   8   :   <   >   @   B   D����   F����   H   J   L����   N   P   R����   T������������   V   X����������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       Y�%Ʉ���>� ۽�R�?nkR�;T���?���?��z��B>�.p>��6�e�p@�R�N��1㠾�, �����Xň@�ý�޾'?�0�Z�N��|�@Z`�
�<��?O��?��"�4�޾��?�Y?�ƒ>|�|?����6z>y�=m�>�@O�_@�]���=l��m�;��3�r>	?�D>"�_<`> �:?;�b?�S�;յ�>�꛽UT=�9e>3#��-�:={�5��+�=�!K�X��<��6=)������؋�=?D���h=�;�>Ճ�n�!���=*�<j�>�3=Ĳٽ���=�m��h�4����=���-���jd>T�;���L       split_indices[$l#L       Y                                                                                                                                                                                                                                                                                                                                 L       
split_type[$U#L       Y                                                                                         L       sum_hessian[$d#L       YC��C[`�C�{C�oBop�B� �B��jC8}A�_�B}KA��A��JBN�s@�Bg��B���A�A�gb@���@�4A�tIA��@rT@@�S�A��A��A�W@�+P?���@kЃBY,�B�)2B(ְ@��@��@@VAT�B@��=?��@͊�?�:
AB|@�Q)@�0@?���@�A@��@$h�A��tA�=@Hp�?�w�@"�A��A�z�B��K?�y�B&o@݂@���?�h�?���?�%C?��?���AB��?�S&?���@jv@���?���Ab�@��@�?�@0"�@��T?�G�@.c@47?�1�@E�F?�[d?�vKA�1�@�i(A���@�(�@BJ�A�1oL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       89L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       ;;��c��PE<� k���ѽ��;�|�>IJ�����@㾥�g�n ��T�<���>�E>��3=nkU��-��e:�=�RO<�ya�ˁI����>H_��R��>B/��ie��,>S`��]��J�=ȓ��Y��p9�>mYT����=�<�>��D�c>�n����F����=��>��-�j\$���W;�>[�W�>g��Y�>� �>�5ӽ$����_�b�>Ϯ;�ꪁ�ӨI>��tL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       ;                              L       idi@L       left_children[$l#L       ;               	      ������������            ����   ����               !   #����   %   '   )   +����   -   /   1����   3   5   7   9����������������������������������������������������������������������������������������L       loss_changes[$d#L       ;@^�? ��?���;�p >"�?gU?��            >Bp�?��?���?N�    >��    ?S.�?�n�?w�O?���?*Ms>���    =�?t?*��?B0�?5X�    ?�%?FȂ?3AW    >��=�}�?��=>�,4                                                                                        L       parents[$l#L       ;���                                               
   
                                                                                                         !   !   "   "   #   #   $   $L       right_children[$l#L       ;               
      ������������            ����   ����                "   $����   &   (   *   ,����   .   0   2����   4   6   8   :����������������������������������������������������������������������������������������L       split_conditions[$d#L       ;��u@?:0?ܭ�@��	\Ϳ#�-�)B>��˽#���|���V?�b?�C�?��>R�*���a�]h>��D>���?���>�q=�f��|侾���B�R>��P?�i��o�g�i>mf#�N�4��"ͽ`�?Z{e?�?�?[�ּk�w=���)6L�,������<���=��н������:�~��W�=(�ߟ=΍�=�s˼E�k�������=�7{�̴���%>I�L       split_indices[$l#L       ;                                                                                                                                                                                                                 L       
split_type[$U#L       ;                                                           L       sum_hessian[$d#L       ;D�A�)(DS�A�4�A�DqB,bAxf�?��?ق�@�piB=�}C�.UB+@�
"@���?��B�{Ap,C��@���@�8�A��?��@|`BA<r�A��AM K@.�C�H4C��@q��?��@"Z?@b{A�E�A(?�^@:T�@YciA�A��A5KZA(��@�w@�eC� AգB��@��?��?��^?� @M�?���@��A:?�T�@��%L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       59L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       %;�<����g��<��!��ؾ=���1[<����AS�T��>�it=2���y�=>_���b������wu?�(<�?G=D�Ծ���4��@��C�<�p/� PO=a2R��H-;�9�=x9J�>3��߂���9�<���۞c>�4Q���L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       %                   L       idiAL       left_children[$l#L       %            ����   	����                  ��������   ������������               !   #������������������������������������������������L       loss_changes[$d#L       %?�:�?�%)?�P?���    ?x    ?�>�>g��?C�>y�`?>��?��        >�[0            ?'�r>��$?���>�]@>�]�>�Bx                                                L       parents[$l#L       %���                                               	   	   
   
                                                      L       right_children[$l#L       %            ����   
����                  ��������   ������������                "   $������������������������������������������������L       split_conditions[$d#L       %?p]�@,�=?��?���8�?�*F��j?B�1��>���?Nv@._.�-��<dr��:־֡���G>0�;�#��!&�\��;�?��,?�����A����<�2�^�:�x�<��-�d=��-��;?����o=��b�L       split_indices[$l#L       %                                                                                                                                      L       
split_type[$U#L       %                                     L       sum_hessian[$d#L       %D*�bD"gB��D!*�@�5�A���A �xD{\@ץ�A�y�@"?`D�
B�*�?�� @�~�A�f�@�L?�!?�_�D q@��RB�/;Aں@�q=A4��A�c�D �R@k�-@I�vBbH�A�+�@�,�A!�c?���@B��@���@��L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       37L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       =����;;����9�j�"=Єܾ�)I����=�s�"�7=�?T>��D��/�>��x�\2>W�[���x�;��<N<8>\)?d�+p�<�J�K�>���0=��R��@$? }��"#=�Y���6�>�ٮ����?:%�>�ܫ���>�^����?���SI�	�>�rþ�#a>;Z)��#(<�5�>Q�������ڞ�>�C9>
�V�[�=/����?�>����A������^�>��V�`L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       =                               L       idiBL       left_children[$l#L       =               	����               ��������                     !   #   %   '   )   +   -   /����   1   3   5   7   9����   ;��������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       =@y6?�>>�*�?�1R?Z#�    ?=�?e��@
�n?�w?2        ?� P?;��>�@?NO�?��?���>?°?��?�8=��?o.6>��">�P?%�a    ?H@2?�u�??;h?���<��     >G:                                                                                                        L       parents[$l#L       =���                                                     	   	   
   
                                                                                                                       "   "L       right_children[$l#L       =               
����               ��������                      "   $   &   (   *   ,   .   0����   2   4   6   8   :����   <��������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       =?:h��%Ʉ?�]׿��@��_?��>:�f��?�4?۹�ԟ�=���=��޾�v=�O��W\����@9�0@^?�|9�S��� g�G� ?��@)�Ľ���>�0?�|?x�.���4?Ü�>�ŵ>_`�?uY?��y�=�%��۔>��30��5h�%`> �����=`Ҙ���;�s�={����H=�,=�P�=&�����<S��Y�=�f�hH������q�=牅���L       split_indices[$l#L       =                                                                                                                                                                                                                             L       
split_type[$U#L       =                                                             L       sum_hessian[$d#L       =C��nC��lAz@NCI�qB�T�A>��@m9yB՚�B��.B�pAR�?�h�?�
jB�vlA��BհBv��B���B	�c@�/@;�B�i�@��A��~@��|A���@��?�HIBpiB��Ad��A��@R�@5L@�m�?�,+?�J�B���@�m
@:�*?�o�@XW�AW/@C׮?�:�A��R?�Yk@@zG@=�wBY�@��9BX�{A.<@���ATjA�5�@jP�?�I`?���@]�?���L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       61L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       M;T���c�<������g��c.;8�=�{����=&@�O��=�׏��c=S��=�n>�>���5>H��`��>wM���>������T�=��>�W����=�[�>هQ��2�=���>�-3�O0.>�r�<y� �u=	X��J�Ƚi$��q>�#�?4n�=n���h>��$���>���>h���-@#>�j�=�-����,>T|~�����ف�<�?#��<����5����%>���Gzξ�˿��<�֔>7v���>�,�>�뗾
苿i[L��/�>�lB�B��=m\>��i�r>��4L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       M                                       L       idiCL       left_children[$l#L       M               	      ��������                        ����      !   #   %   '   )   +   -   /   1   3����������������   5   7   9   ;   =��������   ?   A   C   E����   G����   I   K����������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       M@6�#?q|�?��7>�Ш>�z�?�mI?�oA        >痢>���@G%�?�+h@�>�}@>��R>�p    =���?���?h��?���?��T?�'�?�_:>���>n@>��=��                @ �?��?L�8>��>�@�        ?��j?�.�?=E�?GY    ?�    >�@>���                                                                                                                L       parents[$l#L       M���                                               	   	   
   
                                                                                                         !   !   "   "   #   #   $   $   %   %   (   (   )   )   *   *   +   +   -   -   /   /   0   0L       right_children[$l#L       M               
      ��������                        ����       "   $   &   (   *   ,   .   0   2   4����������������   6   8   :   <   >��������   @   B   D   F����   H����   J   L����������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       M��8\>��l?�VF@pc? P�?����e��1<G�!?7��>T�v?~(P�F�?��>mf#?\�8?��u���=�u{=��|�n�?kj�?�N�0Z�?l�R>^�@*8F���i>�=윤�x�8=҉�;�+���=����G��?K��e!l=���>X��>�8�O���u�<�=خ�?��"�O摿+�ھG�|�>��B�=~�˼������a��>D��;��Z;��_�=?ߌ�o`+�)���6'�;�=[�(�9z^=��=ܴO�&�������b>�[�i��<�C�>���W�=�H�L       split_indices[$l#L       M                                                                                                                                                                                                                                                                                    L       
split_type[$U#L       M                                                                             L       sum_hessian[$d#L       MD�B�ID�2A�3�A�~�C�49B���Az�P?�y|A6��@��AC���Cb��Bk��A�A��@#�?���@��C���A �oA�CY�B6wAV�@���A��4@ع�@�j?�$?�#�@(I�?��B��)C-yp@��h@	"�@��4?���?�(ECW��A�1A��A5u�@C�@��x@ )Ac�_@&�%?�Qx@�e|?�n�?���A�?�B�[4?�C+�Z@ �@s?���?�m@I@�\3C#Z4BR�EA�~�@���A��*@>�D@/�A��@- ?���?�f�ASA�?�>�?�qNL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       77L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       -;��<)�9��0�<��4�F�<����Bx=�����=���f�����;�>�N��\�Ȼ�\.����=
ڨ>�3���:A��~��i.>j�>��x=�=-���>�Γ�٤���i>z<�q==�*i?d8ᾊ��=9��<)\����1>sGҾ�7�=%�>ї�=��rA���a��L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       -                       L       idiDL       left_children[$l#L       -      ����         	                  ����   ����               !����   #   %������������   '   )   +����������������������������������������������������������������L       loss_changes[$d#L       -?��?�d\    ?{��?B?q��?��>��F>�1�?f�?e?p��    <s     ?	Z8>˔T?J�o?R�h?(��    ?EQ�?3V�            =��H>�o�>2Q�                                                                L       parents[$l#L       -���                                                     	   	   
   
                                                                        L       right_children[$l#L       -      ����         
                  ����   ����                "����   $   &������������   (   *   ,����������������������������������������������������������������L       split_conditions[$d#L       -?��?�1<���?ܭ��h�>cV�3�L?�@^���?�C�>��ֿ�J��?	�K��X��S����@�`�?��޿A�咿9穿�=���<ίн�6�@�=�~?��l=7��;�!}<��>��;p<_(;K<����=���ԩa<F�=���=xs��Zž?���`�L       split_indices[$l#L       -                                                                                                                                                                  L       
split_type[$U#L       -                                             L       sum_hessian[$d#L       -D'h
D%�L@���D��A�n�D�IBX�@��A���DҔA���A�1Y@��@D#?�L@�%�A���D��@�kA��@��	A�O�A5Ê?�<�?�Ӌ@aE@��@�D�A/ܠBR�gD tX@]W�?��_A��A�^@�uzAdjA��?��?��m?�1@%��@�~}A�e?���L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       45L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       5�]$�;ؾ����G��=��&����n�:�Z)�]��=|��>��
>�8��ڙ<8#���?�9�O>;�߻�u?(�9>:>�_��&�8������y=�y;Х��%�>�Qh���>�>�l��_���H?1�J�"�>�Vs�g�'>��Ӿ��'��$��;>V->�E]�=���>�(v=W�ھ��e>]����jl>����qWL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       5                           L       idiEL       left_children[$l#L       5               	����               ������������               ����      !   #   %   '   )����   +   -   /   1   3������������������������������������������������������������������������������������L       loss_changes[$d#L       5?�?�2�>�HD?���?5     >��b?,/�?��D?g�?��            ?���?$}@?BX�?��?�`k    ?�;?��q?�K�?1y�>в�>Ͽ+    >�S�?=�?�v?�u�>�7$                                                                                    L       parents[$l#L       5���                                                     	   	   
   
                                                                                                L       right_children[$l#L       5               
����               ������������               ����       "   $   &   (   *����   ,   .   0   2   4������������������������������������������������������������������������������������L       split_conditions[$d#L       5?:h��K�l?�����@��?����?�8;�QB@�ڽ�?L=�׾(��z�Ծ�B?�H�?��?��>J�?�=��p6�>7H0@�@ª?�+���_�>��6����a��@9�0>�Ӭ����n�>U9�Cvx=��$���~=����T�����
jW=����l�=���6	=��<�v���Hz=�
����=������L       split_indices[$l#L       5                                                                                                                                                                                               L       
split_type[$U#L       5                                                     L       sum_hessian[$d#L       5C��RC��5AWÏCC��B���A+�@2C��B/��B��pA�?��P?���@%��CMA�u�A�a�BM�B���@��@��@���C�@�o�A��Aj��@7��AzrcA�a�B+�AA��:@��X?�q�?��"@�t�C1A6��@�׫?�_�A���@@0]@�=AY=@�%A	pQ@.\A��A���A�<�Aն*@)�@tI�?�uL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       53L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       9;/���<~�C���ʼ��-��=`CоIv�>��ȾQx�;�#=��>bF����>�*��E�>�r����e>���=1��-�<��>���=>�`>���>����q��g[=�G�>j�<W���zw�����=�T`=�9��I>�p�= �Y���y=��
>�iS�=U5�W'�>����A��=��F�{��=�p;��/��t��E�>F	��dea>��"=Qxu? ��L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       9                             L       idiFL       left_children[$l#L       9         ����      	                        ������������   ����         !����   #   %��������   '   )   +   -����   /   1   3   5����   7����������������������������������������������������������������������������L       loss_changes[$d#L       9@�5?��8?��C    ?�w?�L]?���>��q>�v�?��=?���?��|?�S�>�            ?I�L    ?P�n?�+?N�}    ?��>��        ?>U�?�d?9c?�P    ?���?��G??<g�    >;�                                                                            L       parents[$l#L       9���                                                     	   	   
   
                                                                                         !   !   "   "   #   #   %   %L       right_children[$l#L       9         ����      
                        ������������   ����          "����   $   &��������   (   *   ,   .����   0   2   4   6����   8����������������������������������������������������������������������������L       split_conditions[$d#L       9�M��?p���������?��->�C,?�վ?Υ��Wm�@=�D���@/1�H�J�;nA=(�3�)�>�m?�~�>�?D��_�����>.��J�?�-=8���n�@�?�{6���n?�#�8,�>� |��>]G�0Zܾ?�X�x�w<H���_=�=��˽c3���=ۍ�hpV<�4T���(=w:�j9�F�3 8=m�3��	�=�4�<{]Z>�cL       split_indices[$l#L       9                                                                                                                                                                                                              L       
split_type[$U#L       9                                                         L       sum_hessian[$d#L       9D�kA�W�D+�AY�A�?C���C�i�@��@9|�BU)CdFcC�K_B �-@�
�?���?��?�9�B�p@
K�C5p�B;WC��@��A���AW�.?�2@E��B� @�[�A�y�C"�J@�+1B(B���C3TA��T?��AG�?�@�A�M@C՚@��@+�-@�6�AIX@Bo�CEhA���A�?:B���A��B���B���A&v�@��?�� A6�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       57L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       /;��q<S��xQx<�c-����`c����<�*��t�p>��'��57>,�f<��T��Ͼ�l8<�su=�|q����=ק��A=c���Q���/�ҁt��w���h>�vp�3�p�T:>�J�����ߴ.=�^#;�P=�44�>�>�%������-�R=�c=?P�ʾ�d�>_��:���'QL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       /                        L       idiGL       left_children[$l#L       /            ����   	            ����   ����                  ��������   !   #��������   %   '   )   +   -��������������������������������������������������������������������L       loss_changes[$d#L       /?�~%?iN�>̒`?MO    >�f�>�8?@�0?9�>�v    >���    ?1�R>-�t>�߸?��=�]�>��        ?2ǚ?]��        >�p�>Ka?5�?\z]9��N                                                                    L       parents[$l#L       /���                                                     	   	                                                                                    L       right_children[$l#L       /            ����   
            ����   ����                   ��������   "   $��������   &   (   *   ,   .��������������������������������������������������������������������L       split_conditions[$d#L       /?�q�?�5^��%�@��������?��?���@5��@
R�=�N����=O:?�վ�����@@�n?�J��-�<3ϖ�َ��ν�0ػرӽ��Y@l�>��P?�Z�@Q�??��=��0���8�<��^;��<���d�#=�`k�=(A�;O�)��<�C�>zt�߫�=�"�9,:�����L       split_indices[$l#L       /                                                                                                                                                                          L       
split_type[$U#L       /                                               L       sum_hessian[$d#L       /D$-xD��A��vD�@���@�'�ASMD0�A�4�@ږR?�E3AC:�?���D֔@�$�A��Afb@B�/@rFv?���A#e�D=�BY��?ν�@r�y@���A?��@���Aj9@�A?���?�@$��CnS�C�Q�A��A�?�@M�f@�݅@~��@c�&?�P�@Ϻ�@B3:?��?��L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       47L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       ;�=��:�3��Ѽ�b!=�H��Nj�C�=T K��j>���=W�[����>���;��>9�s��;��r��bFy>�ʬ��И>�= 񃾫B?!�> ���㞏�:����#�><3.>���>�Ծ�e�=�r=�^>>��z��H1>�����=I>��=K8���� <>�u;fo��.N��0n�Á5>¬<`�`���v>��3�*~���e>�m��h�>0pѾ����>���L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       ;                              L       idiHL       left_children[$l#L       ;               	����               ��������            ����         !   #   %����   '   )   +   -   /����   1   3   5   7   9������������������������������������������������������������������������������������������������L       loss_changes[$d#L       ;?�~2?�P>Ջ?���?H�-    >ܯ�?Z��?���>:x?Q��        ?��?X�>vc�?kp    >��\?$r�>��?ġ�?:��    >��<>�H�>��?=�>�R    ?}�?��?��?��>�|                                                                                                L       parents[$l#L       ;���                                                     	   	   
   
                                                                                                           !   !   "   "L       right_children[$l#L       ;               
����               ��������            ����          "   $   &����   (   *   ,   .   0����   2   4   6   8   :������������������������������������������������������������������������������������������������L       split_conditions[$d#L       ;?:h�?\Kb?�]׿d�>"B��s?��:�zH�I�"�c?ĽP�ս�^�=��P���<�� >�M|@J����>ͻ�?�?���?[/D�� g>BS��I��@������?̗�@!r>��?��nqؾ{�*?���?t�O�^�=��)�#X$<)��=�m�<sݳ���;d�':��N�����=�6;����*�>R�L�־�>
���=S������>��L       split_indices[$l#L       ;                                                                                                                                                                                                                          L       
split_type[$U#L       ;                                                           L       sum_hessian[$d#L       ;C���C��CA<p�Ct��B{R^A�@EWuCD�B�u�Au��B=�m?�%x?͉qB��@BunA�%B��?�
EAe�yA���A�B�EWAOL@2�BF�Ajv�@�}B���AF�@� @״�A(��@��`A��>@�SB��?A
X�@��E@V<�A&<cA�n�AW!?��N@��c@�4B��@��_@�C@�N@�)�@o@�M@�D�@	�V@���A��@E�d?�Q6@�+L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       59L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       7;%Y���	<W�K��K���;�X>{�Ҿ@�=�$<��v��0�=j�Z>݌}��0���S�;��>�g�> �E��E*�CU>4�qjӾ�������<�/>��Y����>��ݾ;I�-W���N=k׾�W�>����ҽ�X����H��쑼�+��s��<�޴�]�1>�7�&XW>������
>��o>��f��>�-k�@k���V�>1�>í���L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       7                            L       idiIL       left_children[$l#L       7         ����      	      ����         ����   ����                  !����   #   %   '   )   +   -   /   1   3��������   5������������������������������������������������������������������������������������L       loss_changes[$d#L       7@ Ao>�i�?A\    >O�?j[�>��=�@    ?��@(>�u     =5��    @D�?�H�?uݪ?�(=��t>Y�    :l� ?=Z?��d?j��?kc�?���?5�L?`ۀ?�J�        >%Y                                                                                    L       parents[$l#L       7���                                               	   	   
   
                                                                                                         !   !L       right_children[$l#L       7         ����      
      ����         ����   ����                   "����   $   &   (   *   ,   .   0   2   4��������   6������������������������������������������������������������������������������������L       split_conditions[$d#L       7���ļ�@�Z��-?v�?�6�>��J?_��<���?���;���5 >��b�2X�G�<n�X?^�?ڈ�UD�>͑��ٲ�/;?bV�^�E�[5{=+־o��x%?"�t�tn<5���ǜl�Xw�����Н��W���4̽�4�<Rl���=��ܾG�6=������>�C=�4��R��P�f焽�h2=;�=��T�3�L       split_indices[$l#L       7                                                                                                                                                                                                   L       
split_type[$U#L       7                                                       L       sum_hessian[$d#L       7DL�A�I D�yA��A�DD	�AI��@ά<?��2C�R�BH+�@݉�@���@�u�@ m"C쁫A�[A�}FA��x@�d@�6a?�&[@;�)A�g�C��3AƁ�@4v�AS�D@���AP
�A��%?�:�?��@f�z?���?�թ?�کA:yv@��4A\JC�@p�A��k?�d�?��?@�ۄA��?�(�@b��A �j@=X�A.uA&{�@%]�?��L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       55L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       #;h�<�ɧ�ǲ<b�?C⽴薾�J�<�p���K׽W���ͼ=+Y���&;���=�ٖ<�]��nb<�N(�8"�?/�4=8�m�=���=�+9��3���O=�'}>��X?z�Q�E->7�=½r���>cI�H=|L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       #                  L       idiJL       left_children[$l#L       #            ����   	      ����   ������������         ����                  !������������������������������������������������L       loss_changes[$d#L       #?�?h��?J*�?9��    ?F�>��?��    ?��            @�)@�H?�N    ?:e�?�<-?�?��]>D��?|�                                                L       parents[$l#L       #���                                               	   	                                                      L       right_children[$l#L       #            ����   
      ����   ������������         ����                   "������������������������������������������������L       split_conditions[$d#L       #?+�?'�>G��@,�=>0��>���R?�^=��'�?�5^�	H><M���?[�p?Ş��R"��QC�o�>��>�^�;�[>��ʝ>�<�3޺��v��^�<�b�=�@�>�T1�ls�=[�7<�#��D�=0݋�pI�L       split_indices[$l#L       #                                                                                                                               L       
split_type[$U#L       #                                   L       sum_hessian[$d#L       #D!S�D/BE&�D��?��qB#HLAy�D��@i�B#9@�(�?���@D��BNt�BAz@N�C�Bf�n@�fxB8�@��A�~CVT%C�f~B,.�Aj��@A-�@�HA���A��?�q�@��%A�_{@�z\L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       35L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       K�(���,=������r��)��=��A;���7�=1d���>_�M�< C>�=��þ]L�>�j��{�����>��k;����b��<���6E�>�s?�b2���k=�����=� i�А=��8�?k��o >7d���>+��>���#���X>�[�>֎q�+�7����<uc=�ze�
�{=}4�?U�>Ibf??X ���>
	�>��'��+N���]�j	>>�i_����=CYr?;?���=t�1>6�O?�ռ��G�c��Ԕ>*�Ͻ�s>����,�=�<���>���L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       K                                      L       idiKL       left_children[$l#L       K               	                        ����      ������������      !   #   %   '   )   +   -   /����������������   1   3   5   7   9   ;   =��������   ?����   A   C   E   G   I������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       K?��)?خN?5&�?�?1�x?~8�?�e�>�pU>9��? x�? �?J�\?7$�    ??��>\Mq            >ި�?0��?�N?"y�?B�?%� ?E�?�`�?o�y                =���?��?[~?/�&?s�?�Z>pJ         >���    ?TP�?0��?��?R�D?&S�                                                                                                            L       parents[$l#L       K���                                                           	   	   
   
                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   )   )   +   +   ,   ,   -   -   .   .   /   /L       right_children[$l#L       K               
                        ����      ������������       "   $   &   (   *   ,   .   0����������������   2   4   6   8   :   <   >��������   @����   B   D   F   H   J������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       K��(��q�1���Q��2迍�t���=�Zx@����(h?���o<��b�c>��?�լ��=�M#��ɻ�1Ҿkx)=Х*@'}�@
�{����AO�=�ľ��G@R���<�f��F���+�D
����R�t�b?�(��_�@ ��>g���F=�ԧ�[l �M�ܿ{2a���0�2l;?;�Z@�>*�<=q�H>e�ͽ�l=%�=�4/��ɽ��׼�k�>rm��YY<jkV>7ಾ�<��=[,>3�ͻ��6�T���=L�,��V�=�h��h�<;Bk;�0�=���L       split_indices[$l#L       K                                                                                                                                                                                                                                                                             L       
split_type[$U#L       K                                                                           L       sum_hessian[$d#L       KC�17B��~CH{/A��+B��3B�y&B�}7@j�aAt�~BA@�B*��Av�#BТ�@�q�B�6@[�?��TAc��?�G�@j�B2��A���A��@QͪAB>�A��B�b&B���@��?�8�?�~�?�@@z�A�&XAh/A�ļ@9�AH<6@_��@��?�N A'<e?��A"�@���BAS�Bp�B�^�@F�?���?�<�AS�;A�a�A��@�dYAb�A�f?��
?�rA8/|?�e�@�r?���@��z@��O@�#n@�J�?�)#@�ZA���A�A���A|�DBp��A L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       75L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       /:�U�����<4�(��6��)B����<�k��	_���ž"��>ʄ<���>�P�=T5��q9��߳��_ľ	��<��=���>���P�_>Ap�u�*=�p�x�={��T��=u�q����>�à>��b<��U��y�m��>���G�ÂP=�F�>�,2���<�Ž�Υ=$�A>�a�>9������L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       /                        L       idiLL       left_children[$l#L       /         ����      	   ����      ����         ��������            ��������      !   #   %   '   )   +   -��������������������������������������������������������������������L       loss_changes[$d#L       /?��.>؈�?;N�    =�Z�?��y??��    >ҭ?l:&    ?�s>t��>xt        ?l��?>�a?"�{>d��        =�:�?59f?��>؈l?�'�?��?x�>���                                                                    L       parents[$l#L       /���                                               	   	                                                                                          L       right_children[$l#L       /         ����      
   ����      ����         ��������            ��������       "   $   &   (   *   ,   .��������������������������������������������������������������������L       split_conditions[$d#L       /��u@?:0��n�և�	\�@S@�Z��q����V�N�8=�۾��0>��J�*���X��9?N��?^�9����@8$>���zhs�i>����ĿB��>���?���5�?��@/�|=���=�l<;H�����>�񺝉z��a<�T�=�Σ�!z�<?�(��<E�=���=_'3����L       split_indices[$l#L       /                                                                                                                                                                       L       
split_type[$U#L       /                                               L       sum_hessian[$d#L       /D�"A��D
�2A�g@�7B?�dC�N?�J@��B/��@~F�C��gA�%@�G�?���@Њ	B��A�]C혡@�X�@��N?��n@]CA��AA�$*A<l�A#��Ck%Cp'@+��?�?�T?�!2A�;A*�G?�(�A���A��@�/A �@
��C3,NB_�5C\.OA��?��?��(L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       47L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       1;[�<E��?{<s`z��}���	꾲ܾ!�q<�\2���=Tg>���?F>uB����>^�G;�w�=��d�k�>E�%��^v�p9����z>�e��qO��D�j0>�&�hǾ���<G��>���%u�GD�
/�>����y�M�>�>��j�d�T���T�'N�<��=���Z����>��> N���R�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       1                         L       idiML       left_children[$l#L       1            ����   	               ����               ��������   ��������������������   !   #   %   '   )   +   -   /����������������������������������������������������������������L       loss_changes[$d#L       1?���?$+I>�x�? `U    ?;ò>��?�6l?�|4?x�?_h�    =��?D.">�# ?�*�?MK�        ?J��                    >ō�?�t?�g�?Ug�?4v?(�3>� �>��                                                                L       parents[$l#L       1���                                                     	   	   
   
                                                                                      L       right_children[$l#L       1            ����   
               ����               ��������    ��������������������   "   $   &   (   *   ,   .   0����������������������������������������������������������������L       split_conditions[$d#L       1?p]�@,�=�'9Ϳ�!&����>�
J��A��oͿ`���l���$�=�O��c}������=�Kj�X �=־NP?~���>(��"��f>	u��Tƿ[l ?yH��'\���i>��@�Z���Ƚ-"R�%��=�>��ґB�v�> xr=�ͳ��:3����H��;�@J���Ӽ��>�=�a����L       split_indices[$l#L       1                                                                                                                                                                               L       
split_type[$U#L       1                                                 L       sum_hessian[$d#L       1D�D1�Aأ�DR/@_��A��AG�A���D�k@���AA�O?��2@��@�-�Am�0B�oD	x�?��E@���A{z@$�R?�@�@��q@HD!?�.�A.a�@}�6A�VA#��@�(�D��@�@\ڽ@��@��*@K?��@e$=A���@u@���@��?�h�D� A q?�-@�K?��#?�VL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       49L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       ;��W;��=��-ݽ ��=�ɝ��L�<�8=�L�2�<�b>7���xK>�"p��ǣ=E����V�"�=�aŽ�8�>r,���l�>�g�<��սMh����?�a�|m=�>��}�\T�=�2�=�R>֛�>���������3u?!����%=S�����>�4��l�=��*���� v>���Q)C=�E�>�">3T�����>�ݥ��	]>�۠��	L?���.�L��� <�g+L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       ;                              L       idiNL       left_children[$l#L       ;               	����               ������������                     !   #   %   '   )����   +   -   /   1   3   5   7����   9������������������������������������������������������������������������������������������������L       loss_changes[$d#L       ;?���?i�J>�pL?�R�?�_    >���?��?�
?6FJ?*            ?�	D>�cp?DL�?�?R�? 9�?i?�?��[?ab�?6>�1H    ?�?[	>���?ic?'6�>���?]�    >��f                                                                                                L       parents[$l#L       ;���                                                     	   	   
   
                                                                                                                 "   "L       right_children[$l#L       ;               
����               ������������                      "   $   &   (   *����   ,   .   0   2   4   6   8����   :������������������������������������������������������������������������������������������������L       split_conditions[$d#L       ;?:h��%Ʉ?�����?ͭ���&?��b����?
G�?Ü�����=�)T��+�zy��cX��W\>�X?�6N�Ƥ�>k�o�|�:c�;��e@6�@>'�ۿ"��sm�?*-ܿN�?�ao=+�?�>0?�_X��p�>A������<~_罞�d=�>����<�����L��[=ז�z�Q=* >r=W2{��=�=-���
=��Z��>\>#�ƽQ���&�;��4L       split_indices[$l#L       ;                                                                                                                                                                                                                      L       
split_type[$U#L       ;                                                           L       sum_hessian[$d#L       ;C��fC��A!*�C4��BݴE@��j@x�B��B��\B�b�B�5?��?��}@�2B¸jAɡ�B_�BBz�A��A��B@���@��XB���@���A�� ?���BZr_Br�AL!PA�RA)�A�+nA'm�?�d@��?��L@��EA��B���@W`?��A��l?��5@vDcBKA�k0A�@�r@��-@�Ah@�C�@��@�z�A,sAvX?Ϻw@+�(?�M�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       59L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       7:˭���9�<+#���ͽ�d:��i>�2�H�z>|����=P=о�>�m]��^=�X�H��>͓S��"���[<�+�>�c�>R��GLo=�4����ݾ��߼޽V>�s�/�=N>�xs�<��E>���t~�>�����-H=�8�պ=���4),>�i3��A�bŚ�H�=�q�>A	 �T\>�O¾��=I�4>�h���QP>�W�>Β�=�� L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       7                            L       idiOL       left_children[$l#L       7         ����      	                  ����   ������������         ����      !��������   #   %   '   )   +   -   /   1   3   5��������������������������������������������������������������������������������L       loss_changes[$d#L       7?�J?@��?1<�    >�?(�>��>�f�>A��?���?5o>�Ky    >�)            >�{�@h�?G    >��F?��v        >ſ�>Դ�>�u�@=�?�L@ �?V�3>��4?�=���                                                                                L       parents[$l#L       7���                                                     	   	   
   
                                                                                               !   !   "   "L       right_children[$l#L       7         ����      
                  ����   ������������         ����       "��������   $   &   (   *   ,   .   0   2   4   6��������������������������������������������������������������������������������L       split_conditions[$d#L       7�M��?p��?ܭ��?�?��-��6�)B>?��W�(�L�,�*@/1�]�>�8�FA=���pŝ=���?7�޿"hj?�^=>o"�9穾��*=	���T�@Ao�>�ŵ�)���#cx>��;�[>�V��@P?���@s�N_<�C5� <i=h��X1i>
ع��[��*�?$=��=g���~�o=͒齦��<q�?>>���a�=��h=��q<�ŚL       split_indices[$l#L       7                                                                                                                                                                                                      L       
split_type[$U#L       7                                                       L       sum_hessian[$d#L       7Dn�A�JD.�AX�A��D FBd�@���@-CxCp��C��0A�K�@k�@p�K?�I?�F0?�@�A�8C^�C�I@es1AiJyAaMG?�K@+��AI@°AX/WCP��CV�BTf@�t@� �@���@��A1�v?�Dx?�
�@�-U@2�`A+�AZT�CB�xB�6�C[�A�lOB/�@X��@r?@y�@�c�@�Q?�=�@#�@nV�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       55L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       #;��<X5x�S<.`�?i���|�˨T<V����+��Ͼ�K�|#��L<��ܽ@<z6����;��=�fQ;Q����TM��w�=�&2=�p���[=A��W�>��Q<�3��'_=�$�>33Ѿ�+�>ySR���L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       #                  L       idiPL       left_children[$l#L       #            ����   	      ����   ������������                        ����   !������������������������������������������������L       loss_changes[$d#L       #?y�%??\�?%C>? �`    ?&ȸ>4p>�I�    >�>            ?h�|?�;�?:^�>:-<?���@��?��?8I8    ?
#�                                                L       parents[$l#L       #���                                               	   	                                                      L       right_children[$l#L       #            ����   
      ����   ������������                         ����   "������������������������������������������������L       split_conditions[$d#L       #?+�?'�>G��@,�=> �>�����>����A�?�m�ƣ�)�*��r<�5��]�?7��?@�u?��?�뺪�!�~��~x��\�?p]�<=����;<g����i�=��;��
���<���=W
���g�=��e�9t�L       split_indices[$l#L       #                                                                                                                                L       
split_type[$U#L       #                                   L       sum_hessian[$d#L       #D4D�B4�)Dr�?�wB��@�snD��@E�^B	��@j�n?��@��hC�4C�A�*@��C�AB��C��A�%@0�Aۆ�?�E�@S CT�KB��nA�)<B�=|B���Bv�|@��A���A��A��SL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       35L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       Y�?��ќ=��W<����0�r>w��=tk='��$7Q��k?���>���>J�����=�t�<��>�n羫�c=��߾�5��+|Ҿ:=�݃�Q�>���-��>�C��ԁx=�9A���n> ����>@=�C>����վ��.�ޙ�>�X)���E�J}���I> ��=�	���2?+�Q��<�j���Gz�,�>��d���Z>U?��={h<�d$�x��>01��O�ܾ���g��M,=:7�=�ܟ���=�`9>��;M ߾�?�� �a>�A�u�>�Dٿ�>�A>́���þN^�>��^=y'c>�ɲ>E66��<�>+�uC[?>�<����>�]����L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       Y                                             L       idiQL       left_children[$l#L       Y               	                                    !   #   %   '   )   +   -��������   /   1��������   3   5   7   9��������   ;   =   ?   A��������   C   E   G   I����   K   M��������   O   Q   S   U   W����������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       Y?n�%?�W�?P�?��?�NW>wh�?��?U�?9�:?x�?	��>���?|>j^>�cf>� =��=��0>�;E>k�?��H?�J�?JB        >Sk_>4�        ?&�C?b]?%�@?�        ;� =�>I <��        >n��?(��?A��?�p    ?�">`_        =�/x?(�?0�O?3j�?�                                                                                                                                        L       parents[$l#L       Y���                                                           	   	   
   
                                                                                                                 #   #   $   $   %   %   &   &   )   )   *   *   +   +   ,   ,   .   .   /   /   2   2   3   3   4   4   5   5   6   6L       right_children[$l#L       Y               
                                     "   $   &   (   *   ,   .��������   0   2��������   4   6   8   :��������   <   >   @   B��������   D   F   H   J����   L   N��������   P   R   T   V   X����������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       Y?\Kb��r2>���>x��>����¾�o?g(?!�ʽ�r+?��@�b&�>��>��`?�"�>~}�Q����]D�Xň>WJ>��?1�?���z��>ט>��O�eΖ���<��@A>?���j׳@*5<��> �j?�~��6C����"�����r���8���F��>*X�@/�>'t��Q�?TTF��-�0�a���п��>BET>(�?�Mp;�ޒ��#/=SnͽyI	�	�7�<$⽨\�<_u�<������=	�>Ur:v�Ya�9�>&[�*�=�k��=�N=.�h��x�w��=�q<�~	=ݾ�=l�u��)=�}g��(j>e����=+k=����L       split_indices[$l#L       Y                                                                                                                                                                                                                                                                                                                                L       
split_type[$U#L       Y                                                                                         L       sum_hessian[$d#L       YC�RSCi�3BsU�C*�*B| %A��5B"߱C�A�qA��QB
2|@�DAE�[@�5B�C[�@�A�@�צAe.�Ab��A��AWs�?�V�@�.x@S0DA�J@7-f?�	AC1A���B�lPB��?�v�@PT�@��;@9]�@���@#��AU
9?�%
@�;�@��	AI�Agm@V*A2�;@ �?�J?��@��@�I @��a@���A��
B�QA��A���@S�@�Հ?��?�Wq?�d@:V?ϸ?��Z?���?��@�ǂ@y��@�u@�u�@�g�@���?���@�:@rDx?�F�?���?Ɓ�@�S?�7y@�{"@h��@-�@3��?�IA��@g;L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       89L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       C9�-|<k�ƾ�zP��((<��>np|�͜G���U��kG>�8�<����j�<!�>ܟ[��+g���>[>��j���t�ׯ�=ߠ�>����>��>&��U��> ����A���5�نQ>#�$���v�q��>!Q+�l)<�c>c���9D>Ъ���t������>�ޭ��S9��2>>�F�>��{��9N����=��<�g���>��6=`tV���g>1� > �|?>@.E�`+�
4�����}�{>�_�Nr>c�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       C                                  L       idiRL       left_children[$l#L       C               	                           ����      ������������   !��������   #   %   '   )   +��������������������   -   /   1   3   5   7   9   ;   =   ?����   A����������������������������������������������������������������������������������������L       loss_changes[$d#L       C?�iQ?��?O>��?&��?�k?
�>:��>��?G>d=n@?��R?�ܣ>�Y�    =��>�J            ?z,^        ?~�?�k?���?�J>"[�                    ?+5�?��>��@?7��?�G�?tФ>&�?<ve?>I\?6m[    >Zp�                                                                                        L       parents[$l#L       C���                                                           	   	   
   
                                                                     !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   ,   ,L       right_children[$l#L       C               
                           ����       ������������   "��������   $   &   (   *   ,��������������������   .   0   2   4   6   8   :   <   >   @����   B����������������������������������������������������������������������������������������L       split_conditions[$d#L       C��n�?�@{6?�a@\~?�^=>�9�?�8V?�!��O8��4?0\�;��>eI>_�?mG���6=�s����K���>��V=-=�G�Zl>��?^�?ڈ���ݽ���
����=DW_���@ +>��?�?#�@?D`�?��?@1�?�b??��ÿtn=�q�;������=�T�=�a���^��c=�;�{�����=�M�<��4��ǯ=UZ'=b>� =f��,�%�л��<��+�=7:�w�=�<�L       split_indices[$l#L       C                                                                                                                                                                                                                                              L       
split_type[$U#L       C                                                                   L       sum_hessian[$d#L       CD
�BJ�C��6A���A�_�C�M�A4�bAe\�@��4A�a?@w�VC��[B#�@��@�ԿA;50@(��?��z@�@o�YA�c?��@��C�4;B��~A2΄A���@���?��yA'K�?�I�?�4E?�	�A9&Ai�A�O�C��>BT��A�v@齈@w� AW��A��C?Ş@22�A ��?�,<A]@�_�Ay�o?�C�9�@�dpA�R_A˩�ATT�@�/@�y@�b�?�P�@�A�y@v
@�8A k?�M?��L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       67L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       7:��O;�㲾W�z<b�?�1�
���Ǿ�MD<�"��c�ʽ�M]�������>����6@��'�<�p>������7c�T�L=��j>@�S�cL�;� ->4�k?�6��<;�ᾅ�پ��><��>�D��V��>Vq����<�Y۾�\8>V����v�?�=�}w>=.��RȾ�BP>N+�ѯƾ����l>���=�f�?Q����Q��b���@�=�J;L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       7                            L       idiSL       left_children[$l#L       7               	               ����   ������������         ����      ����   !   #   %   '����   )   +   -   /   1   3����   5��������������������������������������������������������������������������������L       loss_changes[$d#L       7?W?,>���?�>��*>�xc=���?��?_�>ͨ�    >���            ?|Q>��<?gW�    ?%�P? �    >�$D?��?KR>X�    ?r�n>Ж|>_�p=q�>jt<^6�    >�?4                                                                                L       parents[$l#L       7���                                                           	   	                                                                                                     "   "L       right_children[$l#L       7               
               ����   ������������         ����       ����   "   $   &   (����   *   ,   .   0   2   4����   6��������������������������������������������������������������������������������L       split_conditions[$d#L       7?�q�?g(>�� >&kh> ݼ>�0��=�&W?�n\�VJ<���� �
=�믽����N�)!z=�{>>����!<?��??2k�=gC�����?�Z�>��8�:�B>C��?2v�#=N�A?��?�Y�=-4�>,;�8��"=��-����>3�<�c\=�Ѽ�ɽ��O�=wf�����º�W=���<��>5�?��b�����&�<��GL       split_indices[$l#L       7                                                                                                                                                                                                     L       
split_type[$U#L       7                                                       L       sum_hessian[$d#L       7D�D� A���D�A�)�A%��@��C�B��<Agm>@��DA�B?��|?�P\@�7�C�k@�
�B�0�@�*�Av�@��?���A ��Cۊ|By@�z�?�@B�pqAV@�~!@ߵ@R2�@�?��@�S�C�p@��B�?�w�@�K�?���B�AB)M�AEZ?�-�?� �@�� ?��?��R@c�?��	?��M?���@��-?�a�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       55L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       7�t�a;�Ě��n��٦=�u��A����;V��s�#>���=��E=��͛���I�<�0= w[>�E�<�'>�2�<��K>�6澶���"��U�<��n>k0�c��>�V��O-x>a>�j=�-��� [>�����d�s�=�=w�+>ʉ���������>����M�����>�(O=��ݾ�o�<�=>�R<D���?/��=��+L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       7                            L       idiTL       left_children[$l#L       7               	��������                                    !   #   %   '   )   +����   -   /����������������   1   3   5������������������������������������������������������������������������������������L       loss_changes[$d#L       7?Rw??��=[�?���>��x        ?2��?� >��>�rJ>�v�?c��>>v�?
��>��;cv ?87�?A0>�<8=|�P>�| ?A�E>+�`    >�;V>jZl                ?^�P>�c�?��                                                                                    L       parents[$l#L       7���                                               	   	   
   
                                                                                                           !   !L       right_children[$l#L       7               
��������                                     "   $   &   (   *   ,����   .   0����������������   2   4   6������������������������������������������������������������������������������������L       split_conditions[$d#L       7?�VF?G�?�V>��^����N���L>�zd�?'�?��|?ԼL?g(�0�O@�?�@��V6�f�8?�ݤ?�<����Q��>cz~@5
�>��<Av?s�����=�g�x��=/Du>?�?aP�?�@^@�Խ��W�Ƌ<)"<���=�
ܾ
��=9 ���U=��.ž	Dļ�f_>��<�B=��S";�IO>�e;k=���>S)�<�SL       split_indices[$l#L       7                                                                                                                                                                                                       L       
split_type[$U#L       7                                                       L       sum_hessian[$d#L       7C��C�� @���C`Bdg�@Z?��CIf�A�|@�YBF�nC+B@�<AYy0A~�@;�#@�oB)@�RCK�@wƦANBZ�AH�?���@[P�@�U3?��?��A?�� @\gyBpm@���@�Z?���@�
C�?�<@/��@�ե@7��B'�@ə�@:]�AN[?�*?ُ�?�~j@�2B�*@|+@
`�@��@*>�@g��L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       55L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       79�оO�D</y��s�>00 >���;�K���_=VUY>�*���` >�yN��a'��8I<{�þ�_��׾8�>�����6? �W��9�;�m<(u>b������=�m;뗾��?"�>s�����d��g�=��T<������9<S�J>�?+�h��=>xܦ�R�����6=�ܾ�C��?�3��Q<0|�>\'�=�þl��>V����cL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       7                            L       idiUL       left_children[$l#L       7               	            ��������   ����      ����      ��������         !   #   %   '   )��������������������   +   -   /   1   3   5��������������������������������������������������������������������L       loss_changes[$d#L       7?��_?�9>���? ��>��7>���?
�H>�t<>���        >���    ?{��>�w    >��=H�        =��>���?��>�#�>��=��=�o                    >�0=�à?S�?BN?q��>�i                                                                    L       parents[$l#L       7���                                                                                                                                           !   !   "   "   #   #   $   $   %   %L       right_children[$l#L       7               
            ��������   ����      ����      ��������          "   $   &   (   *��������������������   ,   .   0   2   4   6��������������������������������������������������������������������L       split_conditions[$d#L       7��8\?7�޾���?��P����?e۾�n?U�v���0=� �� ����ǧɾ@V�@{6����� g?��x=��M�4�A�R~�?RP<�O�
?�^=>�9־�#\;�l�:6M齙M,>C0=9V��T����@
�0�B��?���>p��>eI>%�;���5�=�Q1�|���A<8�<���N�j�[>#����;S��=��<�L��4=?4���2�L       split_indices[$l#L       7                                                                                                                                                                                                     L       
split_type[$U#L       7                                                       L       sum_hessian[$d#L       7D~ A��{D��A�>}@;w�@о�D ?A|�@q�?�Oo?��l@�O�?ấB��C쀐A��@��\@*w?�m=?��@e%�AK��A���C�Q�A%��@_�@!?��?�R\@ �?ȡ�@˚�@� �@x��A��:C�"�B!vg@��@��?���@�^?��S?���@�@�(@͠?�0q@"DA�q�C��A�S(A���A�C @���?´�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       55L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       1:�-�= ������<��(>�*�������=
��������7%?\�Yh����)�=���ķx���?Y�>�㼱-�?�J���<��<7�j����>=�i>ҧ�������1�h>���j�g�>��U��[S��K>-�ؽ�7�Sn���V��>�,�{!�=���%�0?Y����y�����?��L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       1                         L       idiVL       left_children[$l#L       1               	����         ����               ������������      ����      !   #   %   '   )��������   +   -��������   /������������������������������������������������������������L       loss_changes[$d#L       1??�K?�mX?�`?Rb?���    ?i,�>���>"    ?E$d@F��?TN?�<�?��            ? ��?y/�    >��?k�?=�?��>$J@?�%j        ?.�?�Xs        >��R                                                            L       parents[$l#L       1���                                                     
   
                                                                                       !   !L       right_children[$l#L       1               
����         ����               ������������      ����       "   $   &   (   *��������   ,   .��������   0������������������������������������������������������������L       split_conditions[$d#L       1�.p��X��V@B�9�C!��5�?��z�R�s@Q�?��u`>w[F?��@+�߿Ss����]��u>���>`���3�>�Y��N�?cF�>ƶ^?����Em�?�@=�ɓ��aC�P$�-��?���о�'������Z=P`���۠�}Q�������9=8uh����=&��Gm>��s���G�˴%>(пL       split_indices[$l#L       1                                                                                                                                                                                 L       
split_type[$U#L       1                                                 L       sum_hessian[$d#L       1D�C�*�C��C�sx@�Ʉ@�C��C�!y@��?��@��C�}�Af
C�\C��@O��?��@Zlx@5��C��?���A��@¨C��@��9@g�C?�?��@��=C��?�t�@�N�@j1h@�B��+A��b@�?��@̺?�+�B�AXB�?�i�@C�{?�%�C�+�?�)�@ �jL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       49L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       9���ҽ���=e(��"� r�_�=��։c���Q��.����;� ]���v>��=��'��|���Y��r/>����>=5��=6k����<�f	=� `��WI�~m�<m�k>�P��nl���V�<�-@>����@�9L=`D>��B>½����s?))���>K?<o���7��+�>�F׾��S>�>W�2�CT.��>�>a�=r}=�[�z�ւ>GTL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       9                             L       idiWL       left_children[$l#L       9               	         ����            ����   ��������         ����   !   #��������   %����   '   )   +   -   /����   1����   3   5   7����������������������������������������������������������������������������L       loss_changes[$d#L       9?D��?��?>�?Oz?!;�?^!	=��    ?&YZ> � ?ח>��    ?T�        ?V{>?���>�H    ?S>�gj        ?-��    ?xyn?{6�?�h�?��&>�ξ    ?�O    ?!�Z>�)?O�                                                                            L       parents[$l#L       9���                                                     	   	   
   
                                                                                       !   !   #   #   $   $   %   %L       right_children[$l#L       9               
         ����            ����   ��������          ����   "   $��������   &����   (   *   ,   .   0����   2����   4   6   8����������������������������������������������������������������������������L       split_conditions[$d#L       9��(�l�1��@��=��L�t���ѿR���~b>�բ?�Y��mQi�=m�>	�?�լ���پ	D;�B�C!��q!<Y��?�T=�^���X�-G>@R��5��!{r��º�ǖ���?s���  ���p"=ۀh?�d�?�������>�[=�U��W>J�ɻ�J�>#{��šv��4e>���Y1=�=����je�
%�=��<�~X���� �t=:U�L       split_indices[$l#L       9                                                                                                                                                                                                          L       
split_type[$U#L       9                                                         L       sum_hessian[$d#L       9C�yHB���C7~�AG�B���B���B���Aw?�t B���A)Bՠ�@k�@�?�B��?�ۢ@�<B^�RA�>A
�\?��iB���A���@!��?���B�:�?�>�A���B�Aq'AU�U@��~@�<:B��#@�%�@��9ApUQB{��@,��?�/�Aq[\?�K_B=�@� ?�13A#��@G��@"�?�xA:��B�T*@��i?��>A#L@��B
�FA��L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       57L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       7:9\L��T�;�&���\��o���w>�d�G𼾓2�;>����6	�� D>J?L�Zc�=�k����<X@�$C=J�F>�HW�1G�=�h>ّ>@�0��n+�I�^=e�p>��x<_�����I P�p.f>��=*x ����>�p��j"���Z]>�Ǿ�,B�f,>R"ؾ��?CI=�z��� =~�D�?.y>�ݕ����w�Q>�9���s>>�fL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       7                            L       idiXL       left_children[$l#L       7         ����      	      ����            ����               ����   !   #����   %����   '   )   +   -����������������   /   1   3   5������������������������������������������������������������������������L       loss_changes[$d#L       7?X�N>�߄?��    =���?$�>��\>3�    ?�n?
��?!n>��    =���?�,?K`$>�Zh>��[    >�^�>�C    >'t#    ?�|?9��=� (>��_                >�[�>�>�/?Cn                                                                        L       parents[$l#L       7���                                               	   	   
   
                                                                                       !   !   "   "   #   #   $   $L       right_children[$l#L       7         ����      
      ����            ����                ����   "   $����   &����   (   *   ,   .����������������   0   2   4   6������������������������������������������������������������������������L       split_conditions[$d#L       7����?:0?ܭ���	���X?�C��T�z�&������#�-�H��h88;�A:���>�|4?�b�!��?��<��=�#�<wͪ�]�>�C�����4��������}�d>��޽[ھq3����=��߿`��?�@^@�+�����
=�#������=N=|)ѽ��F>;��= Q�1hg<��ýej�=�	�w��#�#�z��>�ｿ�$=e'�L       split_indices[$l#L       7                                                                                                                                                                                                       L       
split_type[$U#L       7                                                       L       sum_hessian[$d#L       7D�$A>?KD�'@���@��C��WA�?s@��*?��=C�%�@�$�A�RA��J?��@l|fBJC�%@2�y@M@l
@�>�A�L�@�ִ@*?���A�8ZAC�t@%�OC���?�	2?���?�(D?�q�@h� @I�@�9BA,|�?�H�?���A*�Aq�A8�@]��?�G1?��mC�/PB檇?��H?�@�@ �?���?��H@d�@��@�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       55L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       #:��;��H�ɓ�<+�����<0'>�A3=�M��[�<x�E��*>y{���[�=�����;<5->ʿ��z���_�r�I>�����4A�Ҭ�=w����>�w?.h�E�5=�*�>���=�wU�J`�>@���T���JL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       #                  L       idiYL       left_children[$l#L       #      ����         	����            ��������               ��������         !������������������������������������������������L       loss_changes[$d#L       #?4g;?#,    ?&>É�?c    >�>��^?[�B>�|o        >�3>���>��>��?�	        :� �>Zٶ=�E`                                                L       parents[$l#L       #���                                               	   	   
   
                                                L       right_children[$l#L       #      ����         
����            ��������               ��������          "������������������������������������������������L       split_conditions[$d#L       #?��?�1<���G?�*F�h�?ܭ�>��@	@���?�C��3�L=�����nM=�����@=��$?��޿�J��>ѽ��_>�����ƾ���<�Ƽ��=,J�>P�J�mW�<���=ĲQ<����r�f=3e�7b̾O�L       split_indices[$l#L       #                                                                                                                              L       
split_type[$U#L       #                                   L       sum_hessian[$d#L       #D<�D^b@^v�D9IA��D�T@��@_��A��UD��A�+�@��?��@j߹AV��Dw@@�ZEA�2�@O�H?��@ �-@���@�V�C�z(C>�@U�@?�ĕAc�A+H�?��?��`@b�b@�&@}J@�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       35L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       5�]��;R�@�������y=���Ʊ��ʫs<�$�	�>���=&�C>]�O����f�a=R߷=4�>��<>�>~K�V�i?���}9�>y
���۾��l>�W���!4���4>�	?:z�=��8����<�[�?@�8<�܎���T��?)P=�"=�`3�>&�X�R��]m?$h>�T=�۾��	���=�,(>��n�l�'����>�E�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       5                           L       idiZL       left_children[$l#L       5               	��������                        ��������            !   #   %   '   )   +   -   /   1����   3����������������������������������������������������������������������������������������L       loss_changes[$d#L       5?!�?�<eh ?]�B?�x        ?��?t�5>�?��?�v�?P��?8�N?`i        >���?V�v>G?	>�?L?�a�?"c3?�?n��>�/�??i>�
`?u��    ?���                                                                                        L       parents[$l#L       5���                                               	   	   
   
                                                                                                      L       right_children[$l#L       5               
��������                        ��������             "   $   &   (   *   ,   .   0   2����   4����������������������������������������������������������������������������������������L       split_conditions[$d#L       5?�VF>s4?���g�?� ��o+��4$��'\?�տ�V�@P�Nv4��)޾,�m?D8y<X%�=��?lQ�?�A��[&���Z�Խ�R�;Z����?�����?��?��n>_Ơ�񀽿��<��>g;�;޻�Y2�Μ>J�<��㽆�O=)aແ�2�8>EI�=�2<��Q��8r���&<ڛd>
�v�����j3=�S�L       split_indices[$l#L       5                                                                                                                                                                                              L       
split_type[$U#L       5                                                     L       sum_hessian[$d#L       5C��?C��O@��C-� B�z�@H�e?�RB�BZ�f@��+B��:A<�9B�rB�WA��?��@��)B�A$ɬ@�NS@�b B���A�L?A�CiA��E@���A[��BxP�A�nf?��Avs?���@�ۚ@N[?��rB��@��?�FA�[A+�@�S@��<AXl?ƴ'@=��AqP@� �B#�9A�k<@��AU{<@��u@�arL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       53L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       ):4e��9�<���x��>(�;��>��R����=��>�揽�GS<�D�Ѩ(>�3b=�f���h��h����X>��R;�+>�C<$�@���}m=�B;;�=;�A�X<����e>���<�䛽CҮ����U:	>p�;��>�P>&�ٿ|�=��Q>̆�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       )                     L       idi[L       left_children[$l#L       )               	            ��������      ������������      ����      ��������      !��������   #   %   '��������������������������������������������L       loss_changes[$d#L       )?82
>�V >�>'>���>w�*?'p�=Gx0>��>^;�        ?4t>���            >d�|<�    ?E�j=���        =/��=�i        ?-�?�+U=R�                                            L       parents[$l#L       )���                                                                                                                          L       right_children[$l#L       )               
            ��������      ������������      ����      ��������       "��������   $   &   (��������������������������������������������L       split_conditions[$d#L       )��8\?7��@X�?��P����@Gh^>���?U�v���0=��y�*�@,�=>k�=��C<�᪾	r�� g?� =��c@
�?W�z;E��7�g��#\�fx�:�|��hp�@
�־Xň��`g;��!�j�ѽ�/L��?=��:�J�>
��=G�Ҿ-bq<�
b=�n�L       split_indices[$l#L       )                                                                                                                                                   L       
split_type[$U#L       )                                         L       sum_hessian[$d#L       )DF�A� mC��=A���@3RC��@9�	AZ�@a��?�'-?�xC��i@1"�?���?��0A 0�@�R@�^?��C�Q�@�^�?�b<?��L@O!E@��?�n?��C�&HAt�@�Q�?�2�?�l�?�դ?��f?�nC��+@N@Z��@�z�?��l@��dL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       41L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       /:{��<&6w��jp;��*>��7�:����}�<\,���6e<��c��j= �Ⱦ�Q%<=w>���4��>���=�E��n#k���q��$c>��J��sr<_�Ⱦ��=�[��[J�<L�>�6��H>X�-=X���:�=�Tc>��<�(��	�]��Ň><���ܾ��,<��[�ɶ��P >��ϼ�VS>7hL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       /                        L       idi\L       left_children[$l#L       /            ����   	                  ����   ����            ��������   !����   #����   %   '��������   )   +   -������������������������������������������������������������L       loss_changes[$d#L       /?)�? Ή?�$>�cz    ?'�?7��>袲?4�?�a=�8P?"�    ? (�    ?:�=��B? �B>��b        =1�     >�	�    >�ˁ>�#�        >���>�~<� �                                                            L       parents[$l#L       /���                                                     	   	   
   
                                                                              L       right_children[$l#L       /            ����   
                  ����   ����             ��������   "����   $����   &   (��������   *   ,   .������������������������������������������������������������L       split_conditions[$d#L       /?+�?'潲��?�G�>~!��tB�Ž�?�p�?_O�.$��`�>����?��Q>ˀ��w �����пW�������D?����WV��*���[���>�a��=�A��0>2$>�,n����<�eD=�$�<��%v
�� <=�$Z��iս�_;�����r�y�=�Ƽ�e=B}L       split_indices[$l#L       /                                                                                                                                                                         L       
split_type[$U#L       /                                               L       sum_hessian[$d#L       /DSfD
�B$JID	��?�1WA�nIA0L�DՃA���A�o�@���@��_@���D�-?���A��_@'[�A��@�l�?��#@o�C@�$?Ӌ3D/j?��M@�	NA{.?�,�?̊�@��KASȷ@a�@Uw�?�C�?�ށC�-C
c�?��@j��@��5A(c}@��?��?�sTA:�L?�ž?���L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       47L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       3�p?�;R���A����E=a�n�������c��y�=�>���<[l�"XE�ǡ�����>*>��Mh�>ǂ��zX;
�q>�����S�> �:��6/��Х>�9p�b�a�j�>Ўн��=a�8?	��>Ig�{��>E~[��A�=���T�=>��8=�!^��t�=gᾦ���(��>�� m�>�a>�\i<��>�U۽`ǡL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       3                          L       idi]L       left_children[$l#L       3               	��������                                 ����   !����   #   %����   '����   )   +����   -   /����   1������������������������������������������������������������������������L       loss_changes[$d#L       3?�>�7K<�9�?D�6>ԉb        ?��>���>� >�7�?��?P��=���?=��?sCi>��}=��    >�o�    >�Ҩ?##�    >Φ    >$6�>�[�    ?4�U>��C    >+�                                                                        L       parents[$l#L       3���                                               	   	   
   
                                                                                                  L       right_children[$l#L       3               
��������                                  ����   "����   $   &����   (����   *   ,����   .   0����   2������������������������������������������������������������������������L       split_conditions[$d#L       3?�VF�K�l?��v>G�@��.?��O�>z�?s�����?۹>�@ �?�~�?�@��?��?\Kb@^��>7H0=���@�?�����3�r>�D���>��6=�D�?v����>%)�?@1»��=l����<���y}=��<��q���H<|����i�JN�=,dV�@��=٧�=��;��=�3Լ��.L       split_indices[$l#L       3                                                                                                                                                                                       L       
split_type[$U#L       3                                                   L       sum_hessian[$d#L       3C�v�C���@v4�C$B��$@4%I?�^C�gAgi�B�~t@���C�A�fsA31@�mYA���B��}@�]c?�vRB���@AiAH-+@�?v@�ʥ@7{?�X@��SAP hAgNA�HB>��@	6�@[�7B��A7aA��@%�9@&9�@dED?��d?���?Ȫj@H�r@�n�@֒*AĄ<@�^@� B(rw@kB?�1�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       51L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       /:�X���<LCt�Ȯ?�8Ѿ��<��̾�{���+��]>�,7�f�^>w�?��<eߐ��L��y�=�|>�؞���"=��>Ѧ��2�2<$F>�.��Vv?=�:�������4�p�>�Iw����<Sg����r>�z��H*<��}��n�=��-���@>>p7�ʢ����>��.<�1>�e�=��L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       /                        L       idi^L       left_children[$l#L       /               	      ��������            ����   ����   ��������      ��������      !   #   %   '������������   )   +����   -������������������������������������������������L       loss_changes[$d#L       /?+�H?Zo�>�ye>"_X?;i>�??�-�        ?!�D<\�@>ڠ�>��e    >���    ?��        >�J�>�        >�l>it>���>��>���            ;�B@?'+K    =ҋ�                                                L       parents[$l#L       /���                                               	   	   
   
                                                                                   "   "L       right_children[$l#L       /               
      ��������            ����   ����   ��������      ��������       "   $   &   (������������   *   ,����   .������������������������������������������������L       split_conditions[$d#L       /��n��R��^�E?�a@\~<�l޿X��-��7�O8��2j�>ܙ>��j>9��@�Z�ǁ>�U�<��=�7%�w��>���=��ĽVEp�Rd��\�X??�v�a��?__��S��u=���?U�F�E�μ�d#�N� �Ӊ�;�]c���=Y轫lM=d����(ѽl�=׍;*�> 	�<8s�L       split_indices[$l#L       /                                                                                                                                                                         L       
split_type[$U#L       /                                               L       sum_hessian[$d#L       /D�B.�C�y�@���BF�Ae��C�K3@�+?��{B ��@[�TA>�M@�@�XC�A�@g�HA�+�?�x�@EA�~@C<?���?�^UC�3�@�zxA)gA�x @��W@��?�5�?�P�@:p�C�?�U�@��@��@�ۑ?�cA���@S�h?��?�?��@��C�l#@u��?�(�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       47L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       59{��;�����<Qj���꽎�ξ�LG<�9̽�db��;E�� ݾ���=�x����G��S�<6�>��ᾚ�ܼ�=�8��C>41`��g�=��,�k��<��]���0��u2?"�Y<�%	��<�?�����G>�ཽ���<��Ⱦ�þ�C3=�����9>��^?t��>�p��j�{>�T�=���?j��=��o�b��{�>л->�X��,	L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       5                           L       idi_L       left_children[$l#L       5               	            ��������         ����            ��������   !������������   #   %   '   )   +����   -   /   1   3������������������������������������������������������������������������L       loss_changes[$d#L       5?��>��>��t>��*=uϸ?��=Ŧ`?��%??B�        >�H�?�)=責    ?d�?��??1{z?�        >�N	            >���>g�X>Ʉ�>���?3��    >�t?]��>S>L>iIu                                                                        L       parents[$l#L       5���                                                                                                                                                       !   !   "   "L       right_children[$l#L       5               
            ��������         ����             ��������   "������������   $   &   (   *   ,����   .   0   2   4������������������������������������������������������������������������L       split_conditions[$d#L       5?p]�?���'9�?΄���>�
J?QN?�{?묬��ຽ��׿l���$�=��%� ��?��L?e�m�)
3?�ۑ<򩸾�\?~����<�h���t&@,�=?��<���?�1ƿ"(��$V��Z�?��D?�/V���;��W������P�<��p����=�zq>���=�!3���>2�<��>���<�����+��#c=�z7=(ٝ��4�L       split_indices[$l#L       5                                                                                                                                                                                              L       
split_type[$U#L       5                                                     L       sum_hessian[$d#L       5DI�D��A�v�D��@y�Av��@̥�D IBE��?��v@!Ǽ@�B�A%y�@3x�@e�kC�R@�2A"�BR}?��y@f�A
-�?�\�?�s�?�~jC��@�qB@T`@@��@+@Ė@�0B��@�aj@/��C��n@[@�{2?��A@�?���?�#S@P�z@9o7?�w�?��?�?�A�N�A���?�E@���?�Ay?���L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       53L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       9�%,�=[��
q�=w�?"�}�M'�;��E�>�Ъ��@�>S����<�G!<Xn�M��Q��>�L�>~T���i>Ö�pԿ�k�TW�>n���=2uɾ�e>�?�ź���Ҧ�/�=̮�>�R*>��U�fｂD�=L��<N�Q>�������<���?��>W�־�O�>S������nҽ����抽y>�ʾ�5�>`�>N ���_4>��h<�+L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       9                             L       idi`L       left_children[$l#L       9            ����   	                        ��������   ����      ������������   !   #   %   '   )   +   -   /��������   1   3   5   7��������������������������������������������������������������������������������L       loss_changes[$d#L       9>��i?�w�?���?:��    ?���?���?B]�?��? &�>��>�X?
?H�s        ?H��    >���=yP            ?�m>�R+?�>e��=� ? �~>�>�P        >�$|>��5>ϓy?k�                                                                                L       parents[$l#L       9���                                                     	   	   
   
                                                                                       !   !   "   "   #   #   $   $L       right_children[$l#L       9            ����   
                        ��������   ����       ������������   "   $   &   (   *   ,   .   0��������   2   4   6   8��������������������������������������������������������������������������������L       split_conditions[$d#L       9�1㠿4�J�I�"?��>Cv0?�R�*��? �}�g��+ͪ�Cu <�������A0��:]A�{Ǎ���=��d=�O���ƽ(�e�#0�~ϱ?�̺%Ʉ>c��=:�?�A���@����V�<��I>d��L��?h���TA��`;x[�=����NB;��>3�==�a����=}��	@X�4������W ��w�>ۭ����=��M=wZa�٥r=�J<L       split_indices[$l#L       9                                                                                                                                                                                                             L       
split_type[$U#L       9                                                         L       sum_hessian[$d#L       9C��B�� C+]B��n@=A�OC��B��WA?`�A�m�@�y�@�0�C	fMB��B?�E8?���A%��?�A�m�@8�?���@I�d?�@A4YB�AyB�U@���@�6�@0-
AD7�A<�m?��|?�H�Ab�@/�DBf�B���B��w@��@��?�<�@�v@5�4?��|?܂�A3��?�0�AX�?�V�?�A�@�u�?�S�?�\�@�N�BU#D@NG�B���L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       57L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       :y)(�Z�S;�\���T׼��*;�E�>�ta�=�>xL:�ė>����p>󆼞�'>�S�;�۾�@A>�*�=l��=��`��l:3d&>��?;��K� Y;�<׾�'H=��I>ؾxL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L                      L       idiaL       left_children[$l#L                ����      	����               ������������      ����������������      ������������������������L       loss_changes[$d#L       ? |�>�L>˻A    >Ǔ�>���    >~�E=�R>�/=9e0>��Y            >���>M@�                ? �Y=���                        L       parents[$l#L       ���                                               	   	   
   
                              L       right_children[$l#L                ����      
����               ������������      ����������������      ������������������������L       split_conditions[$d#L       �M��?p��@7��́?��-@X��=Ǿ�?Υ��(�L@Gh^>��n�FA= �Ի�Wb=�18@,�=>k�=�fK<��<�m��\�@
�?j��:�|����:�I��/$=__>�L       split_indices[$l#L                                                                                                                 L       
split_type[$U#L                                    L       sum_hessian[$d#L       Dp�AD|sC���@��g@�jC�K�@9M@���@�xC��@<L{@`x�?�]j?�^�?��OC�x�@-*~?�Z�?�>u?���@��C�z
@���?��*?���C�@�3@�g�?��L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       29L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       59���=a��\K<�d�>�0��}μ��;��u>	띾���?DҼ9���vf�<��\��� >`HT�328?LHw=��b����?l�E��;1=��= ,��]c5�[����8>��7�j���.�s��>�⏾D�Ϸr�JҬ��6Y���>�s����<'I>S9���iսC� >��ٽ�(�>b`��N���#=��??C�t�������?��L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       5                           L       idibL       left_children[$l#L       5               	����         ����                     ����      !����   #   %   '   )��������   +��������   -��������   /   1��������   3������������������������������������������������������������L       loss_changes[$d#L       5?ϼ?���?uh�>�ǔ?yI�    ?/�z?��^?Y63    ?($d@	�M?C�?P��>H��>��>!��    >[��?@�z    >
� ?D��?Z�?	x�        >���        >�{�        ?ި?��        >��
                                                            L       parents[$l#L       5���                                                     
   
                                                                                       !   !   "   "   %   %L       right_children[$l#L       5               
����         ����                     ����       "����   $   &   (   *��������   ,��������   .��������   0   2��������   4������������������������������������������������������������L       split_conditions[$d#L       5�.p��X��V��Rb�C!��-c�?��z��% '��+l>w[F?��@+��@$4��*��@��p�>u#ÿ)��3�>��]�N�?cF�%`�@,4p����(�?r�Z�,���k��mX=�vF�Q��9��-�� ��h���'��a;./%=}xq�
?��k,'=�8��c�=��m��+D�?�*<�L>k���f\��2>t�L       split_indices[$l#L       5                                                                                                                                                                                                 L       
split_type[$U#L       5                                                     L       sum_hessian[$d#L       5D��C�~�C�ԱC�y@��@�C���CjA�&�?�L@�z�C�W�AJ��Ce��@��A���@�?�@J�"@0?�C���?�+@�	�@��CXr�AS-?��@EչA�~�@��?�:@�1?��|?��0@},PC��Z?ք@�h�@`s�@kxC@�`A�Q @�?A�nA��@,3�?�ZB@<�@��?���?�D�C�
?đ�?�VKL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       53L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       3�?��; F۾�j*<�W۽�{&��9彠Gi�_�>���#�>0���g=�a>Wأ��v��
�B�D��&�>��~;�	t���?��=�羐>�NY��1�>��k�!��콐>��ƾ R>.����rs? ~<=����i>��Q��33���>����y>��<������羯��>O�0�6Y=�d[����>�%�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       3                          L       idicL       left_children[$l#L       3               	��������                                    !   #   %����   '����   )   +����   -��������   /   1����������������������������������������������������������������������������L       loss_changes[$d#L       3>���>��<�P>�A?�\        ?e
?#o9>�2>��>�%?+�l?,&?�$>\��?>�]P>(e�>��|?��    >���    >���=d`�    ?C�X        >3�F=wj                                                                            L       parents[$l#L       3���                                               	   	   
   
                                                                                                L       right_children[$l#L       3               
��������                                     "   $   &����   (����   *   ,����   .��������   0   2����������������������������������������������������������������������������L       split_conditions[$d#L       3?�VF>��^?�
?���?�B���Ez��U�?!�T?J*>̵�?�=;=>d?)X�.�=�(?�A>�H1>��@!U?%%�>�8�>9|�>�y���7��o��,��=�X�?=���W>�D?�&B?.�K���W>1<-��1�=Ѝ���=q�ŏ;=(�G���=��;̣6����	Ѿ�Ҳ�=ymm�Zo8= 	��rO=���L       split_indices[$l#L       3                                                                                                                                                                                        L       
split_type[$U#L       3                                                   L       sum_hessian[$d#L       3C���C���@\��C`�:B�@1n?��CD�HA�G�AΉ�@�'C z�B�aA���@��6AJAR�@���@(Z�B�9B�K?�|wB~?���A�e�@�M�?��A)@O�V?���A?��@/�@$q?�qA?�D]B��@D@AkФAɦDAҎ�AX	A���@�7�@ؿ@�+@�8�@J2A��@��?�{�?�~.L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       51L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       7:�gn�-(�;�j��l��>݄>g�;�Mf���.=E;">�B���=>�T���b�ȉ�<K���B��I���W>w:�`��>��޾�#�:t������=$s-�|=���?�=��������O���&>A�<�#1�Z<��J>2�׽P4����>W���I+�Y�v>9Yw=˯ᾁ��>�l���>��:�!O�&�Z>�4�=9�役�d=3>�RyL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       7                            L       ididL       left_children[$l#L       7               	            ��������   ����      ����   ������������            !   #   %   '������������   )   +   -   /   1   3   5������������������������������������������������������������������������L       loss_changes[$d#L       7?5>��>��W>���>f��>�1>���>���>'W�        >�b    ?C)�>��^    >@��            >P��>��>�[�?aU?~E=� =�(V            >_?	@8>�Z�?7�5?K:?'�?\�                                                                        L       parents[$l#L       7���                                                                                                                                                 !   !   "   "   #   #   $   $L       right_children[$l#L       7               
            ��������   ����      ����   ������������             "   $   &   (������������   *   ,   .   0   2   4   6������������������������������������������������������������������������L       split_conditions[$d#L       7��8\?7�޾���?��P����?fǾ�n?U�v���0=�O��4���8��^�@Vۼ�������� g��h=�V�����>AA�?RP<��a⾆5�?�վ��#\;�l�>?��<ſ/�z�?�۾ݑ�?&1o��ZX?��?A�ڿH�J�y�����B=�k��$�����=^k\<�l�����>	!�5��=���9��ƽHA�=�?a<^��޿E<6��=�b�L       split_indices[$l#L       7                                                                                                                                                                                                   L       
split_type[$U#L       7                                                       L       sum_hessian[$d#L       7D ��A���C�esAo�E@/�@�Q�C�D+A=@Kp�?��?��@�ǎ?�)�B.�C�~R@͙+@�m?��x?���?���@O9�A*��A�4CP�qCvG3@A�u@�?�?���@� �@� �Ax�HAe!C��BL3�C\GA���?��?��?�>r?���@��?�"�@�KA_�@�X@��@�b�C�nBB��@=�C9r�BS5A�:JA��L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       55L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       9��<;,ް��D�;����8<�d�xĽx*s���G<r�g��}{�6���<:C�>��z�u�i��p�=2G������e��'Y<�C��	�/=��?9۾,�=�E>�!��(�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L                      L       idieL       left_children[$l#L             ����         	   ��������                     ����   ��������������������������������������������L       loss_changes[$d#L       >�V�>�5P    >�R-=]�`>���>�@~        ?i�>��X>V.`=b� >�:�>"�>��    >��?                                            L       parents[$l#L       ���                                         	   	   
   
                                    L       right_children[$l#L             ����         
   ��������                     ����   ��������������������������������������������L       split_conditions[$d#L       ?��?���߅�?�P����?ܭ�?����E�ܚ�?�C��3�L?3�ʼ�e ?�?��޿�J��d@,�Y���y��=��bk<(��%�=�>>x��Np�<S=9䎽���L       split_indices[$l#L                                                                                                                  L       
split_type[$U#L                                    L       sum_hessian[$d#L       Dj�Dƻ@#�?D�~@k=�D��AOs�?�da@�aD�A���A��@���D��@���A���@);w@�2X?���?�%@1�C�3�C*@N��?���AQT9A%��@��?��L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       29L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       5��,��`�<<�q ���n����Qr@=��Ⱦűƽ�(�>���.�);�����+t>�d�=@�m>�k=�����=7]<��Q0���0n>�о���=�V�<��:��=��_���m<Gf�>�K�=���ƃ��Ù��&�>!I;��$>��ཁN�������>��;��<�˝��ޅ>�|�=��[��oS>w��>��3=$r�=����JL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       5                           L       idifL       left_children[$l#L       5               	      ��������            ����   ��������               !��������   #   %   '   )����   +   -   /������������   1   3����������������������������������������������������������������L       loss_changes[$d#L       5>ץ�?-Xn>��"=�i�>�T>�6�?oN        =i >���>�>���    ?"�        ?p�?n>�Q�?�=�1�        >�u?0�?}>�PL    >��;=6�>���            >���>�j=                                                                L       parents[$l#L       5���                                               	   	   
   
                                                                                             #   #   $   $L       right_children[$l#L       5               
      ��������            ����   ��������                "��������   $   &   (   *����   ,   .   0������������   2   4����������������������������������������������������������������L       split_conditions[$d#L       5��8�l��?H��!ٺ�3�ؿ i��;���d`�+�u>
+u>�=*�p><X�*�.>	�<�s���r>G�?��=+ֽ��8=4�ǽ�p�>� ۿR�8?<,�?���ƿP?�o�@�F?(,t�C�����7�Q�?,��=�ڧ��+K��C���@=�x+:�N�<Ž���=���<�ס����=��u=�r�<EV�=m�����L       split_indices[$l#L       5                                                                                                                                                                                             L       
split_type[$U#L       5                                                     L       sum_hessian[$d#L       5C��B���C$�q@��B��B�I�B��4@���?��@|�B��*B�']@�%@�HIB~�_?�$m?��Bc�sA�S�B�ġA�@�R�?�J>?��/Bw�A놞A�&HA���@`B��I@^��@�ֽ@p��@@{�?�R�A��@B7�@�JlA�4A]F�A[�@���A���B��s@:�@�?��?�	k@A��A/A^HRA��A���L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       53L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       =:i,���6<K?l�m8=n\�>�f�<�+������>
���h�n>�&5=,H|�rC�<o)n�22� �n�ˌ��B#q>hm���B��=��꾩��>�萺X�=�=���UP=1�4����>�ff>9M�G{=ȉ��ֵ>���Ԥ<+򡾈IJ=��+�J����>z��˧�>�ݭ�0��>Ц�>��7��4Ѿ���>�ӿ<=���<��ս���@�w�ҡ��>L�ཱྀf�>��L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       =                               L       idigL       left_children[$l#L       =               	                  ��������      ������������            !����   #����   %   '����   )   +   -   /   1������������   3   5   7   9   ;��������������������������������������������������������������������������������L       loss_changes[$d#L       =>�4z?��$>��?2E�?HX<=�&L?�U<�@?�&?/IG>Ѕ        ?G�>�GI            ?T�?#�>��>��z    ><    ?��?;��    >Ѥ�?��l?��>R�>�av            >���?'#?�α?s��>���                                                                                L       parents[$l#L       =���                                                           	   	   
   
                                                                                         $   $   %   %   &   &   '   '   (   (L       right_children[$l#L       =               
                  ��������      ������������             "����   $����   &   (����   *   ,   .   0   2������������   4   6   8   :   <��������������������������������������������������������������������������������L       split_conditions[$d#L       =� 5D?I�ҽ!=���E�?ݙֽ�o|��n�if��8����D;��>�<N�b@��>��w�"<<�IQ��B9�Խ�P"?�*��,��=~�����=���=�3�@�4�ٙ�?����H^L�f{�=���?�ڌ<�G��m=!?J�=qZ>b��@>�Ӭ��=���b�=�pj�S��=�a�=� C��?b��U=]ʾH
<��4<뀼�8ݾgü1c(�7	�=u�t��H8=2m�L       split_indices[$l#L       =                                                                                                                                                                                                                            L       
split_type[$U#L       =                                                             L       sum_hessian[$d#L       =C�oB}��C޻�A��B�@H4�C�+@��:A��A�K@ԛ�@z�?�t[AyC��U?��@�*@�wA��A���@��@�_�?��1@��s?�f�C�
�B���@\�DAh��@�:tAL.P@]a@�7h?���@i��?��@˛�C�MAW�`B�Y�A��Ad�@��K@Y�|@b�m?�7�A9Q?��m?�'V@P�L?�	@�1�?���C��B1p�@f��A�A�/�B8�@�pA?�.�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       61L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       =9?R�;��0��[�;�/�>���������C>E=��=�5��m<�o���D<-b���)k>�Y�=¾P��>���a?U>�r�>�+m���6;�n�>�����b��=�/�?�r=�]��R�
Fྒ�B���B>�:��E\��&�<4╾���?�̾�b�=р+��J�	���&c�Ck<>K?d?BSZ<�"���t>~y���4�Д�C��>r�?z�<�����6v>)���%!����L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       =                               L       idihL       left_children[$l#L       =            ����   	                  ����                  !   #������������   %   '   )   +   -   /   1   3��������   5   7   9   ;������������������������������������������������������������������������������������������������L       loss_changes[$d#L       =>��m?/j>���>�t=    ?]�?��?C��?]'e?@�K?M}�? �_    ?�5?{n�>��?���=��t?D>��            ?q�p?G��?��?��=l��?NJ?��>�$        =�H�>�a�?��;��                                                                                                 L       parents[$l#L       =���                                                     	   	   
   
                                                                                                   !   !   "   "   #   #   $   $L       right_children[$l#L       =            ����   
                  ����                   "   $������������   &   (   *   ,   .   0   2   4��������   6   8   :   <������������������������������������������������������������������������������������������������L       split_conditions[$d#L       =?+�?'潲��?�^=>n ��$�Ž�?[�p?Ş��R"���C>����v?Q ����2>��?Fu��H�>}t�>�N>	�<=����Ŵ�?K��>�*��o��?f~���?#;�[>�L���%�dP�p0.�� g>}Y�uv;Y�
�4>|�����<�f��"�&�%]�����j��=s�>i0�;�]*���7=�����4���LK�k�='V�>2-;����Χ�=K�ڽF(ɾ��L       split_indices[$l#L       =                                                                                                                                                                                                                          L       
split_type[$U#L       =                                                             L       sum_hessian[$d#L       =DJDB`ED�6?㶃A�y�A�!C��B<uA9R�A�Е@m>G@�{ C�Y=BI�b@�l�B$��@v��@�Q�Ap:�?�1�@+�?�$�C��N@�{�@�		B+�A@�t@m0�BPG@��?���@2�@.8@�5�AKL@��YC�?�@]��@mK�?�V�?��G@��8@=�-B �?��:?���@/�?��A]�A��@X"�@mP�?ִ�?���@n'�?��0@L�Z@�K�?�X�@�IL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       61L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       �e�>��p����=��+>��B���8;�]ʾ��)��n}>�U �oQ�=>�"2�j�:�7>_'��<L>�:����R�D�;,̍L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L                  L       idiiL       left_children[$l#L                ��������      	��������      ������������         ����������������L       loss_changes[$d#L       >�pd<g@?c�`        >���?>��        <�� ?)K�            ?/�C?U?�                L       parents[$l#L       ���                                   	   	   
   
                  L       right_children[$l#L                ��������      
��������      ������������         ����������������L       split_conditions[$d#L       �p��<ߠ(�o�|=�M=�߃;�l�m帾�滾0���l��=<!>���-���Z�z�c6=����+0�k5:O[�L       split_indices[$l#L                                                                                     L       
split_type[$U#L                            L       sum_hessian[$d#L       C}X�@@d�CzW?��?��r@�z�Ct�G@�%�?�T�@��Cp*�?��W@I�?�n�Cn�AMl�Ca�6@�P�@��OAx0\CRL0L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       21L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       %����Gy�;��߾��=��Y��<�h�ĳ<$鹽�A�>U���tWi=��?�B;�.m=����2�=�a߽����ӟ��J�>������tE<�c�Tsd>�!���Ͻ���>��\;��Y���u>�}�
�g>��?���<5o@L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       %                   L       idijL       left_children[$l#L       %               	            ��������      ����   ��������������������   ��������         ������������   !   #������������������������L       loss_changes[$d#L       %>�K=>���>���>��=���>��G?XA]>���=&v        >w:�>��!    >��                    >�`m        9J8 >��z>��            >&Q�>�es                        L       parents[$l#L       %���                                                                                                              L       right_children[$l#L       %               
            ��������      ����   ��������������������   ��������          ������������   "   $������������������������L       split_conditions[$d#L       %�M��?��Ϳ^֚?sB���潫�e�X��\�|?��$��q=�a�>��P���>$0��Rd�<����=��ܻ۽�ʿ?AhB=�׽6Bp?U�F�E�ξ� g=�W[���_�f5���0�#�-��+Z=f��&7I=��7-q;Y��L       split_indices[$l#L       %                                                                                                                                    L       
split_type[$U#L       %                                     L       sum_hessian[$d#L       %C��uA(/8C�\�@���@#�Ae8YC�38@���@�?���?�xLA(C�@s�r@�vC�.?���@��?��?�Q@���@��V?�D@ �n@0��C��,@��?�f|?���?���@��MC��@|�u?�[�?��k@Y�eA���C� �L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       37L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       79�Ki<�����D0<�m�>�B�������<�V�������?͛���g'#;�+|>hϋ>D�����?A�=ߕ-��8�?FB`�Ԍ=W�<��(���V>��=)��>�&�����>ah->�~x�����'c��o���������>��I��x��� �=��̾�+t�r�O���?��>�f{�%&�=���>�G�8lܿS����������H�>��XL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       7                            L       idikL       left_children[$l#L       7               	����         ����                     ����      !����   #   %   '   )   +   -   /����   1������������   3������������   5��������������������������������������������������������������������L       loss_changes[$d#L       7>�Hr?kAd?M�>���?DOx    ?�R?��Z?�`�    ?$?�:�?!:�?() ?}k�?�Y?!�h    >>/�?:;    >��?&VG>��s>�PN?_Y�?@��=�)�    >`�            ? Mf            >��                                                                    L       parents[$l#L       7���                                                     
   
                                                                                                   !   !   %   %L       right_children[$l#L       7               
����         ����                     ����       "����   $   &   (   *   ,   .   0����   2������������   4������������   6��������������������������������������������������������������������L       split_conditions[$d#L       7�.p��X��V�Un�3�r�!�R?��z�&0�ux��J�>w[F?��@+�߿,6�>W�?�Wy��Y
>h�7�)�?�T*>m�A�N�?cF�>.��?�	��*~�� ��=�k���� �p=�>�=��Ľ�
�3��������꾓'�ґ(��'<�()����c� P=>1cw=�GǽF.�=$�>v+�]Oo�1���G(���`��#�>�5L       split_indices[$l#L       7                                                                                                                                                                                                        L       
split_type[$U#L       7                                                       L       sum_hessian[$d#L       7DZ�C�xC��<C���@ҡ-@	�C��,Csa�Ace�?���@��wC��A:�C[��A��@��A�@@6��@,��C��V?ϲ@�6�@��MCSH�A�eA$#AW�@�1+?���@��W?��?�&�?��MC�'@l��?�ɳ@��O@Y�e?�gC�oB���@��@��"@ ��A��@��h@��@	�@u:@hO�@�ґ@k1]C�=�?�]�?�g+L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       55L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       =��H�==����a�<�Ϙ?U�I69�Ӭn�85�>g�/��1�=%T]���Z<*0�='9�Z��JϨ>��p�ڔ��1>P�S���վ�|��^K�<������>��ϻ%B���B=��>�����о S��b��iC<�>:<�>��1;W>)���5L�E����p? ��<�2���E�q����l=�>�2?�X>@=����x>7N(>�`�����>�>�=v2<s�:��>�o�}�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       =                               L       idilL       left_children[$l#L       =            ����   	                           ����         !   #������������   %   '   )   +   -   /   1   3������������   5����   7   9   ;����������������������������������������������������������������������������������������L       loss_changes[$d#L       =>��}?Y��?BTs?H�    ?;�>?9�?d�>��>bݘ?o�=�@0>�`�?F��?^�]    ?&;=��`>y��=��            >�B_=� ?5�?�+>ք$?74�=�V0>�j�            >؉�    =L�>��?`6                                                                                        L       parents[$l#L       =���                                                     	   	   
   
                                                                                                   "   "   $   $   %   %   &   &L       right_children[$l#L       =            ����   
                           ����          "   $������������   &   (   *   ,   .   0   2   4������������   6����   8   :   <����������������������������������������������������������������������������������������L       split_conditions[$d#L       =�1㠿4�J���?��>)�R?#�+�GϬ�g�=�O?@1�>���@9�0�|sԿ2l;�s_���������"�[�UL���3�J���`�?�C?����ܿ@��kyl�p�?�A����( d��7��K����;aR>�6�?��n?�t��ُ��ܼ�>@��<Q�������<�9������> ��>*�=f�ɽ��*=[�d=������=��<���;�C#����=����ADL       split_indices[$l#L       =                                                                                                                                                                                                                             L       
split_type[$U#L       =                                                             L       sum_hessian[$d#L       =C|J�B�r(C!�B��@�.A�hCrB��A0�mA^#�A�!@V �C��B�+�A&2�?�c�AF�A�@��@@��@��@%3?��C�9@9�x@�TBw�	@�;�@�)*@�B�@6��?�D@�.�?�>@n\�?�LZ@�;�B��AL�?�c�?�wl@+��@<��Bc�@�S�?֖{@u,�@(L�@�@�� @�?���?�w	@�?���@)�]?��B�b�@u_.A��@CmKL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       61L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       !:!�X�QD;����h��>�~;&��U�L���<%<v?_�����;�6>��J�����=��X>PO;H�{;�?>O��>4��Ǚ>��j��vĽ��h<!��Ngb>؉q�����8��BC�<]��L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       !                 L       idimL       left_children[$l#L       !         ����      	   ����   ��������         ����   ����      ����������������   ����      ������������������������L       loss_changes[$d#L       !>�%�=��x>���    =\Y�>S{~>�m    >5L�        >W��>��<��    :�V     >zd>>�7�                >r`�    ?/^>���                        L       parents[$l#L       !���                                                                                                  L       right_children[$l#L       !         ����      
   ����   ��������         ����   ����      ����������������   ����       ������������������������L       split_conditions[$d#L       !��u@?:0�ց��ӱ!�&��?v���8\��&��CV;FH�>?�?73/������ g�sf?7��<��?fǾ�n;%�=x}�������k�(�Ǝ��@V۾���w�C>���J��]r��i5;�.KL       split_indices[$l#L       !                                                                                                                      L       
split_type[$U#L       !                                 L       sum_hessian[$d#L       !C�Y-A�C� �@7I�@�rA@"8�C�_?�z�@�S�?���?�y@�_�C�R�@v�?�`v@t��?�l�@Ö�C�D�?��?��@2�=?��@�4�?�>B ��C�$�?�52@L�]A��A�)�@�9CڔkL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       33L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       =��gz;�Κ���<���U좽|ws����<l�>�^=�
r��x�<������m<\��#?	E���辑�!>yE���R�n���v�>��,:��>	?����>�%H��>Φh>��?�s��>w�վ���=<_e���{�j�9=��Z<M����@�>�4���7�-����x����*�ս�Cx>�]���=g��=S�>��f=�����ŵ>���	?}<G����4�<�wﾺE�>�W��|�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       =                               L       idinL       left_children[$l#L       =               	   ����               ����      ��������            !   #����   %   '   )����   +����   -   /   1   3   5   7   9   ;������������������������������������������������������������������������������������������������L       loss_changes[$d#L       =>��e>��>�-�?�b?A��>wL�    ?.��>���?��Y?wFW?�/    ?��?�-s        ?��F?7s<?Z�0?4�:>f�t    ?	#?��>R�    >� �    ?�V>G�L=R�`?Um ?r3O>��>@�6>�4�                                                                                                L       parents[$l#L       =���                                                     	   	   
   
                                                                                                     !   !   "   "   #   #   $   $L       right_children[$l#L       =               
   ����               ����      ��������             "   $����   &   (   *����   ,����   .   0   2   4   6   8   :   <������������������������������������������������������������������������������������������������L       split_conditions[$d#L       =?
�>"��> ݼ=�&W���=6����͙=�4�=�{>>�n?{S>�V	��ꃽ)!z�;�p>" ����6{?��L��=o�d�]�g>ǁ� ?�?��Q?s�D=��W��	�=���V пcX�U�l>�]Z>7�@?%���9��rI;v����=�q���CܾP����;Ľ9�?�M	 �߄*>k��	D<��<�=��{<��*���@=�p�$��;o�j��;��S�߆�=������L       split_indices[$l#L       =                                                                                                                                                                                                                                 L       
split_type[$U#L       =                                                             L       sum_hessian[$d#L       =D�rD�#AwӕC�kB��nAB\�@U�C��@���A��zB��A�|@#(RC�P�@��-@���?�tq@ʧA��A«�B+�CAě?�oC�S�B�@g�1?�>S@�iC?��AEˮ@���@ˢA�2CB,@�qR@��r@���C���A�tA�%_AaK�@'K.?��@%�P@&�7?�(�A)��?�<�@��L?�@n?�V�@��A���@ʊ�A鵋@9�@���?�*>@ �@:�?�bL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       61L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       ?�?��U�<������3�Ğ�r�
=��S�dT����>9L+�N%�;I(����(>��[=n��>U1��y�*��0��P?<4�>�����w��<��<���M;9�=�鏾�=;>������<A�t���=�,<�"=[�f�+�پ��B<�f�=A�>��i�$�c>��B��\���:>�ܐ߾�>���=K�>�~�(�}�D�>E)��v8=�侽�5ľ�S�>A�����<N�y>�l	>��=��XL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       ?                                L       idioL       left_children[$l#L       ?               	                        ����   ����������������   ����      !   #   %��������   '����   )   +����   -   /   1   3   5   7   9   ;   =����������������������������������������������������������������������������������������L       loss_changes[$d#L       ?>���?�>ӯ�>��2>�V�>��?p�>t�<�_�>���>��>Ʀ>R�`    >ә^                ?N�u    >�h>��v>���>�Z�        >�@E    >9��<옠    <))�?F��?T��?jYM>J�*=r�0>V1?��>]\                                                                                        L       parents[$l#L       ?���                                                           	   	   
   
                                                                             !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (L       right_children[$l#L       ?               
                        ����   ����������������   ����       "   $   &��������   (����   *   ,����   .   0   2   4   6   8   :   <   >����������������������������������������������������������������������������������������L       split_conditions[$d#L       ?��8��q�1��������Ǿ�à�d��]�?��P����G����(z�>N?��=՗�����l����^p>���G?:���*?�r$?Ky���F�:^�?ci\��|��k��$A�;h�%�`}�i��1㠾�V�@*�>:��?���@-�V6�E��=�M��
�e��y�V���K��wN<t��=��N�JH0�*� =l�W���U<�~��@���12=h���;�6;x8+=�?>s#<���L       split_indices[$l#L       ?                                                                                                                                                                                                                                  L       
split_type[$U#L       ?                                                               L       sum_hessian[$d#L       ?CxF�B��CA�@B���B�9�Bo��@,�$@�EnA�B��B��@��@�;HB_u+?���?�_w@���?�vF@���@:�@�u�B�f�B�K�AE@[D�?���BYk?��@oԱ@�?�4w@s�>A�9B:��B��A
 )@��@��BH�m@���?�=@@&6?��?�Us?��@2N�AS�A22@�<�B(�B4P�Aߌ�@ױ�?�:@ A�@���@$NY@%��B9�@}�@ �?�~]L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       63L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       !:d��C$;��H������>�&�;'��9�<���>�2K=��V����;��d��@�=w�x>.̾�����p<1z���=3���	�=�+:�c>K5��P5��A>��+�:��	}>G��>�	����L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       !                 L       idipL       left_children[$l#L       !         ����      	         ��������      ������������������������                  ��������������������������������L       loss_changes[$d#L       !>� �=��>���    =WU�<L �>���>.a[=���        >3A�>p�t                        ?8'/?k�=�L�?�:�?WZ�?*��                                L       parents[$l#L       !���                                                                                                  L       right_children[$l#L       !         ����      
         ��������      ������������������������                   ��������������������������������L       split_conditions[$d#L       !��n?:0�ց���s�>k�->!lž�8\>R,Խ�6=�<[<��>��>��޽��Y<��H=P�\�>�ҽ��!;T���g�$�*A+>�k��[���%C>v�l���s�(�=���`+��$�n=os�=��>��L       split_indices[$l#L       !                                                                                                                       L       
split_type[$U#L       !                                 L       sum_hessian[$d#L       !C��BA	[�C�Sc@.�@���@�EC�9�@P�@&��?�+�?���@���C��u?�Ӵ?��X?���?�W�@:�?�@eC���CŠ@�ScC��WB���A��@�z�?�b�@�{�C�hBը�A��A��$A$(L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       33L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       9:�<;̾���=��!��th��R���PG��w�>�r���;*��>&�@��6����>���>ט.�#Gt���*���>iEʻԂ>�� ���7��&���Z�<�����*>�/�Vb�>��C=��2>[�m���>�J^��=���;��7>�t����=տv�'���#�'�?H�=��O�Sb�>���>�<�V�����	�>�����
0��r>sL�>Y���L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       9                             L       idiqL       left_children[$l#L       9               	   ����                           ����   ����   !   #������������   %   '   )��������   +   -��������   /����   1   3   5   7������������������������������������������������������������������������L       loss_changes[$d#L       9>ü >��_>��Y?�af?>�>�Fp    ?*��?2˂>��?�i>'H�>�jF?)��>Q�8>n�P    >ؙ�    >��>� m            >���>�E�>�g~        >>��>�!�        >PF�    @PK?�b>Z�Q?i�1                                                                        L       parents[$l#L       9���                                                     	   	   
   
                                                                                 !   !   #   #   $   $   %   %   &   &L       right_children[$l#L       9               
   ����                           ����    ����   "   $������������   &   (   *��������   ,   .��������   0����   2   4   6   8������������������������������������������������������������������������L       split_conditions[$d#L       9>]R�`�>��ֿs�C�Vix�X����-#>�V=�+�>���K���ۃ��QB���,��w�מݽC�Y�� g�'��?��J�g�D=�Z��C������@<lgA=Q!>黀��;�l�5�$=�����*?
�
�%,�h��c'�?@1�>�� = ?��1��
��<�@>)�w=�0�}��=�(x=�l��t�����=�_;��r��8�V=���=��]��vL       split_indices[$l#L       9                                                                                                                                                                                                              L       
split_type[$U#L       9                                                         L       sum_hessian[$d#L       9D&�D	 Aó�B++UC���A��/@>�IA��AT��@�^�C�@_��A��[Aɺ�@�g�A5n�?��@�ї?�3�A�)C�<z@��?��>@X#�Ai��A�
�@��k@6��?�9A�@�?��@\�@�ѳ?�Z~AȾ�Cఋ@���A�VA?�@�)@�$@+7�@�ŧ?�=�?�[�?��
@�$?��_A�d�?՟�Agt�C�t�?���@}�A@~>�@��?L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       57L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       A��Do�� =5Bn�ɪξ=�b<��>i!���s:��8��~j=J?�=<ך�e�G>��=7O>��G�o$e�wL��?�>�0<�N�<�U>I�a=	�ؾ�Us>j����;z�>�����>cT��&4>\��6:�+l���>�=��|=HJ�n��V�D>��<>��Q�k�=�'>��'��f�>�:?�j;��������3�Ǽ�A>���}Ͼ�ʾ�Ij�}\`<���?��=��ľ�ME>CŎ��&>�����N�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       A                                 L       idirL       left_children[$l#L       A               	      ����               ����               !����   #   %   '   )����   +����   -   /   1   3   5������������   7����   9   ;   =   ?������������������������������������������������������������������������������������������������L       loss_changes[$d#L       A>�u1?�>>��`>��C? �>���>�yZ    ?��>�0$?(E>�c(>�]u    >ԥ�>���?��>ό�=�    >g��?	�??m�n>�2u    =���    =�Ͽ>�J*?2��>�m<��@            =h    ?y�z>��>荃? P                                                                                                L       parents[$l#L       A���                                                     	   	   
   
                                                                                                         #   #   %   %   &   &   '   '   (   (L       right_children[$l#L       A               
      ����               ����                "����   $   &   (   *����   ,����   .   0   2   4   6������������   8����   :   <   >   @������������������������������������������������������������������������������������������������L       split_conditions[$d#L       A�%Ʉ>z�@���@	��?�U�@�ڽ���z�Ծ��D@=�?��?���>k?�j��ke�>~|��pv@<��>�@P/�?9�>?X<h������?�>Խ��	=��S�`/ƿ2&-���>+D�=���
 ��M�����Z=��?
斾o��?K/�?�6(=�Db���<-�b=̙ɽ�?=0B�>>mL:̟��5�Wr#�
'=������~&�ًM��:;�L>$F�= �C��)�=j��g�>�ɽ�L       split_indices[$l#L       A                                                                                                                                                                                                                                             L       
split_type[$U#L       A                                                                 L       sum_hessian[$d#L       ACs�C�B��C�VA�:�B��B@ܝ�?��PB���AS��@��B�@R@�^�@w�@�a�@�d�B� �@��A�[?�h@�HB��A2��@@��@3@CX�?���@(��@N5XB�>�A�@7RZ@
O�@�"]?��e@9�?��B���@���@P�/@�0�?��S?ʷ:?��?C?�gs?��h@	��?�AiA*�BЙ�@2��@ľ�?���?�/?�t?���Bx�@8��?۫~@��?���@:N@��?��L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       65L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       )9� ��-��;�q边����:��>�̬=�.O����=Q���IU���>���<�)�?	E޾��;$�9>��s�SL=�nZ��w=�L�?L��&�=z�\>���>�>Ϯ��;G>]�����m��>�	}�≿-4�>��4��>�U	�i�Q��)\;>�`L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       )                     L       idisL       left_children[$l#L       )         ����      	����   ����         ����            ����         ��������   !   #   %   '��������������������������������������������������������L       loss_changes[$d#L       )>�2�>��>�8�    >��h>��d    >5��    ?�?��>�[    ?+��>���?bg�?ʩ    >�w>?�V�?E��        ?J�?.%	?('�?��                                                        L       parents[$l#L       )���                                         	   	   
   
                                                                        L       right_children[$l#L       )         ����      
����   ����         ����            ����          ��������   "   $   &   (��������������������������������������������������������L       split_conditions[$d#L       )�M��?p��@7���"W?���R�s=���?Υ������Ss�L���7KC=��+>�F�?���>�Ӭ�J�=�㾿��_?�7?��=	��>t��O��?�Z�� g�P|�=.�8���=���s����=��0�0C�O��>:h�X�\>3��a1���o:d�AL       split_indices[$l#L       )                                                                                                                                                       L       
split_type[$U#L       )                                         L       sum_hessian[$d#L       )C��:Aq�C��@Qug@�(�C��@&R�@��?�:?B��C���@k��?�,�B�)@p\�A��9C�S�?��p@)G�B�\�A��v?���?��^A7�@�0�@��C���?��A?��B.OB��Ao@K�@���@�m?�1@s�@�Xu?���@��WC�@�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       41L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       9F�;v����8�[:>��t;�ԁ�%�u>��=}��<G���jL�M�L��u>�~`;����b�>)��Z@=�6��_<��=��I�W�n>ܷ����=����:>l�پ� pL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L                      L       iditL       left_children[$l#L             ����         	   ��������         ��������               ����������������������������������������L       loss_changes[$d#L       >��>��C    >ѡ=���>���>��,        >�)�>�R�>�m�        >�|$>��?b�>�#>�
�                                        L       parents[$l#L       ���                                         	   	   
   
                                    L       right_children[$l#L             ����         
   ��������         ��������               ����������������������������������������L       split_conditions[$d#L       ?��?�*F��E�?p]�?Nv>cV>���>s<�L��� ">��>��v��YC=�dt�R�s�Yq`>�X��q.?~��4�r;ҙ�=�����B>m׽���<����B�=��齝Z L       split_indices[$l#L                                                                                                                   L       
split_type[$U#L                                    L       sum_hessian[$d#L       D	�:D	J�@PD�	@�D9(Ab�-?���?��C�>�A�;A)�R@e7k?�xC�(A�U�@G)�@�3�@� �B�C�Y�@p�Axo�?�MS?�6@r�@�@�.t?�ɇL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       29L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       1��%z<O�ܽ�}�;�#>��Y�#��=�\�ϧ�=��ʽ�܌��������>�:�;���I6�>���cc¾`�l;�p־^[V>(�&>�S�<'��`�>��>Ii���	><�<��Xb��qf���>��w���۽9e澖��>��ͽ$O����=�?�>��{<�)���$>0��z9[>_}���D[>/���I��=s(EL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       1                         L       idiuL       left_children[$l#L       1            ����   	            ����               ����         !   #��������   %   '����   )   +����   -��������   /����������������������������������������������������������������L       loss_changes[$d#L       1>�;K>�i+>�k>���    >e�t><�<>�F>Ĝ�>���    >���>��>�V;>�V�>�g�    >5:�>���<�<0=��        >��>5v�    >ئ�>�t:    >�]y        >54                                                                L       parents[$l#L       1���                                                     	   	                                                                                            L       right_children[$l#L       1            ����   
            ����               ����          "   $��������   &   (����   *   ,����   .��������   0����������������������������������������������������������������L       split_conditions[$d#L       1>��^>��?�wQ?���=��k>��?�>?Ԑ�@X��>̵���kM?��?��?��Ⱦ���?�R��o?�A>�z��[�>�ŵ>��;IsH?h͆>���=q��@#��.���6�?=����i�=�j�>*X�^zH����=�f��E,s���n=��>J<���=SUk��"j=�!���=Rъ�rb<���L       split_indices[$l#L       1                                                                                                                                                                                 L       
split_type[$U#L       1                                                 L       sum_hessian[$d#L       1Cpl�CR *A�e�CP�?�I�A��A@�R+C6��A��KA��/@G��@�O@"QC,LA$��A�bf@�$A��A"��@�@'��?��/?��tC(�@Y�?�5�A	�A���?�H�@�K@\�?��sA�z?��0?���?�ʄ?��zC��A�.�?�j?��1@��V?���?�W�A��_@�p�@3��@�1�@��)L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       49L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       A:��H��AU=�A�?��;�W?h<��ڿ4!��I�>�@������>¨:�� ����� ��?.,p��,�<<�%<Y����R=z>�R>t:N�EIE���=��ܾ���>��?=���?ot �ޘ�=�W�?>��;���wx>'K>�1���&>ƴW� �x<���?Fǿ�;BzA����e�<TN��ݡ�>�!�?��m���n�&�߻�UH=��<�d��0:f>������'>V��Ogy���=�n�=��>�RWL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       A                                 L       idivL       left_children[$l#L       A               	����   ����                                 !   #����   %   '   )   +   -����   /��������   1   3��������   5   7   9   ;   =   ?����������������������������������������������������������������������������������������������������L       loss_changes[$d#L       A>��z?�qN?��z?���?W�    ? �_    ?ު?��?�)R?��>�@�?�	">o�d?�?;9>�@x?�eV?��    ?0 E>��?!�S?l=�>{h    >-�
        >���=���        >��?&c~?4Կ>�3�?= �@                                                                                                    L       parents[$l#L       A���                                               	   	   
   
                                                                                                         "   "   #   #   $   $   %   %   &   &   '   'L       right_children[$l#L       A               
����   ����                                  "   $����   &   (   *   ,   .����   0��������   2   4��������   6   8   :   <   >   @����������������������������������������������������������������������������������������������������L       split_conditions[$d#L       A>ϛ�>++�>�P���g�D>;���ʾ�(�.$��j���`2��p�>�җ>�ܠ>��p�OXȽX�@�4�^��?vn˾��>eI@Q!���8�?n1�?m{�<�)��k�=��<���iH>��<�ϝ>e)�>:f�?�J?�?�?��h<��3�"W��R�;��>+wt:i_��
�ż�z;~�Ծ��=��1>��P�T��HT?�
3,=\A;�xֽSyH=ŵ8��Mb=��C�xⒾC�=-<��7> ��L       split_indices[$l#L       A                                                                                                                                                                                                                                           L       
split_type[$U#L       A                                                                 L       sum_hessian[$d#L       AC�H�C�5yC.&�B�2C���@(�C,/@�:+A�;�A��C��kC�A���A�{o@��@�8�@�`�A1\�C���C�:?��ZA�hDA	YA�MA> �@ԓN?��z@X#�?��p?֮`@'j�A-:?�{K?��KC�o�B��A�yYA~��@x��@�9?�a�@��u@bXI@_�A-�@��?�O?��p@@k?�V?�&@�8@xxCg�NA��GB�AjA�b�A#z@��oAbX?䫴@
��?��.?��h@ȏ�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       65L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       ����:��Z��=���[�>�v�;rx���>ڤ�=g�=<%^ؽ�gŽN����;���>��}��}���Ir�%m�>%<7"��-(�E��>�߱� ��C�>���X]s��*�;�@~>��Z�-6L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L                       L       idiwL       left_children[$l#L             ����         	   ��������         ����                  ������������������������������������������������L       loss_changes[$d#L       >�1�>�(    >�}	=�;�>~F8>�L        ?=�?fND>yF�    ?2w�?X�P=��?\�8>pw�>��3                                                L       parents[$l#L       ���                                         	   	   
   
                                          L       right_children[$l#L             ����         
   ��������         ����                  ������������������������������������������������L       split_conditions[$d#L       ?��?�*F�Ȱv?p]�?Nv?�J�>���>/�<��?� ?묬�1����?��L?py�"(�?�ۑ>��v<�:@;1�ý�id�mw>�7��$�jb>�c��Ѭ��3K:���=˒�O�L       split_indices[$l#L                                                                                                                       L       
split_type[$U#L                                      L       sum_hessian[$d#L       D	5�D��?�cD8	@�D��AW�y?��?�A�C���B(��A$�]@LDnC�T?A)w�@�6�B�@�9Y@zj�C��@喯@��F@��n@A �@Gl�@"�"B��@��@{��@��?�i�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       31L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       =�u�=�U�
f��˦9>���Jü��L<�V��:?r�=خ<������Gr��=I�m;g��>���䇊=A�r�� }>�ݾ����l�>u��<Ů<�.پ��	>��;�*��zm��{�-�>�i[=�Hh>����<?t>�W?�M��sN>�"ۼf!�>O�;;�Q�>��9��N?�=��ȬN�]�=�Lh���=�� ��]�����=k��>�H߽�.�>PF>�ҽ�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       =                               L       idixL       left_children[$l#L       =               	            ����   ��������                  ����   !   #   %   '   )   +����   -����   /������������   1����   3��������   5����   7   9   ;������������������������������������������������������������������������L       loss_changes[$d#L       =>�<>�v�>�w�?;yl>�s�=2\�>��B?}">���    >�ͼ        >��Y>a��>��7>�l ;r ?=    >���>n<�?uЏ>G�h>��~>��\    >�A<    >5-�            >�:    >���        >�Z    =���>��c>�3{                                                                        L       parents[$l#L       =���                                                           
   
                                                                                       !   !   #   #   &   &   (   (   )   )   *   *L       right_children[$l#L       =               
            ����   ��������                   ����   "   $   &   (   *   ,����   .����   0������������   2����   4��������   6����   8   :   <������������������������������������������������������������������������L       split_conditions[$d#L       =�d�:�zH�+ݩ�����v�C?\Kb?[/D�� g>�ܾ� ���|��و�=��E���?JN;�񃀽�Q��!���c�.$�@'�>�4�h?՜�?#�/��r�`�D�L�ӿC��.�����X=�~n�KB=�s����D=?��>.���e����?�Y�?��@uK:���=⎫����>"�<5E����Ž���=a���� fm�ͣ���It<�_4>+����=y�>	K?�:$ L       split_indices[$l#L       =                                                                                                                                                                                                                             L       
split_type[$U#L       =                                                             L       sum_hessian[$d#L       =Cm��B��B��B�V�A��@��JB��B�J3@��#?�)�A�F ?�c�@s<�B�|�B8��B�&q@�<(@��)@2K�?�nWA�A���BU��@�SB'0-B�n�?��3@��p?���@:��?�&�?��?���A�Q�@�4�A��q?�5�?�{LBO�?���@S+aB̜@��B��M?��?��o@b)?�P�?�"@.�A�L@�e^A�O@|#[B?M�?��@
�vA�̆@�2�@6q�@o�oL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       61L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       9:ŉ����<E��ve�=	yܾ�B<^�~��R]>O�>�����
��]F�G�>��<-8о�Dž=��=� >�ϫ>T��q�Y��	�=!⼾�i$��Ȩ�%�>D��;�(�>]�ʾ�1l=����,��>���=.��ÐT��0;=��>�#D���<[q��B{�ы�>��>�R�����>��[��)r��R>����!�>Ū�>3 v�p��;�tL>�6>b�΀4L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       9                             L       idiyL       left_children[$l#L       9               	                        ����   ����   ��������      !����������������   #   %   '   )   +   -   /   1������������   3��������   5����   7������������������������������������������������������������L       loss_changes[$d#L       9>�?8Q>��?$J?F�>2��?�w>n�p<��?  >�&y=���>�i�    >�~    >�9�        >��d>M&                >� >�OU>�Tq>�:�=���>^n�?X	J>��h            =k�d        >��    >֥|                                                            L       parents[$l#L       9���                                                           	   	   
   
                                                                                         $   $   '   '   )   )L       right_children[$l#L       9               
                        ����   ����   ��������       "����������������   $   &   (   *   ,   .   0   2������������   4��������   6����   8������������������������������������������������������������L       split_conditions[$d#L       9�ǮO?_��^�E@`?ݙ�?U�v�X��4l����\��@/?b��(A>A@�����?&y<$@ =�_�?��?�?��Ҙ<BCI��J�������=�J@��7N���?��?Ja|�M�$<5k��2��m�o��>���>�$@C���.�?qy=�9~�|8��e�=�4��1����=�ǹ��[�=�3#=V�����5;�a=�@�=������L       split_indices[$l#L       9                                                                                                                                                                                                              L       
split_type[$U#L       9                                                         L       sum_hessian[$d#L       9C�;B�oC��NA�hA�uvA5D�C�7&A^r�@��A��n@�"@pʯ@�$�?��YC�I9@�zA5�?��	?�iAd�x@َ@J�??��	@'R�?��"@��n@RqC���@�@�p�@W��@��-A#a?��o?��@��@8f?�]9?�G�C��?��@S�@�j[?���@�
�?�}�@��@�P@U
?�.BA��?꡾?�*uC�]�?��|?�_R?�G�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       57L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       �s0U:U�龙h;簾��(:�J>�k;��ɾ[">�8=]�;"�>~pC�8�f�c;����	}>�[K�<�U�oH=�L�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L                  L       idizL       left_children[$l#L             ����   ����      	      ��������         ����������������������������L       loss_changes[$d#L       >��r>{L>    >��    >��k=WO>b�>��        ?��>:CW>B��                            L       parents[$l#L       ���                                                              L       right_children[$l#L             ����   ����      
      ��������         ����������������������������L       split_conditions[$d#L       @,�=?�4���v?�*F��&�?p]�?Nv@Q�?>���=�O<�"�@B��@SR��1���f�:�M=��c>i��b� �2$=��L       split_indices[$l#L                                                                                    L       
split_type[$U#L                            L       sum_hessian[$d#L       DL�D��@
��D]�?�!vD�@	�&D�AJ?�Cx?�
�D��@+#�A� @/VD4)@I�?�N�?��'@�1@q��L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       21L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       �R��;fƮ��l>���a��=�	�>������<���hٽ�>���9��w>�\�>F˜�L��<S�ƾ>���>뾦x�>s��:0�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L                   L       idi{L       left_children[$l#L             ����      ��������   	   ��������      ����         ������������������������L       loss_changes[$d#L       >���>��     ;�]�?6Qx        >6�?(�        ;*� ?o7    >��?:�?�                        L       parents[$l#L       ���                                                                    L       right_children[$l#L             ����      ��������   
   ��������      ����         ������������������������L       split_conditions[$d#L       ?�VF�p����X�<ߠ(�o�|=ғ=Ѡ�;�l�m帾r�8���Ȱ�aD@>�"�+'P�|��������=�r�=�����=�4�9SFL       split_indices[$l#L                                                                                            L       
split_type[$U#L                              L       sum_hessian[$d#L       Cj�Cg��@"@3�Cd�j?ս?�b@�$�C_�E@Z��?ׅU@�PIC[L�?��6@G��ABǕCO I?���?��j@V�AD]A��CEdlL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       23L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       A:������"<2��
E>��=o�z���!�ҬV����=��>��N='7?�Ͼ[h�;�du>�Q����=��۽�$v?C#�><;��#�=�X��<�m>�Y�=j���ԛ�o�����(>�q��;<>P�G�����>]�Ծ�����K>V��>��<7QO�?��=دX=���=j?�|�"����E����>����`꾠�>fۨ���5�ݽ�X�>�f������>�E1��>~߮?KI'���<<��L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       A                                 L       idi|L       left_children[$l#L       A               	      ����   ��������                        ��������   !   #   %   '������������   )   +   -   /   1   3   5   7����   9   ;   =   ?������������������������������������������������������������������������������������������������L       loss_changes[$d#L       A>���>��&>��>�Y�;� ?�gX?Q˂    >��=        ?�e>|�@?/�>�
<��>�C�?�m�?�x�        ?$?E?�K�?�_x            >��?�F'@@b?M%�?�U6?C�>$��>��}    ?\p5?h>ŉx?)�O                                                                                                L       parents[$l#L       A���                                                                                                                                                             !   !   "   "   #   #   %   %   &   &   '   '   (   (L       right_children[$l#L       A               
      ����   ��������                         ��������   "   $   &   (������������   *   ,   .   0   2   4   6   8����   :   <   >   @������������������������������������������������������������������������������������������������L       split_conditions[$d#L       A��n@\~�R�s�N�c�4�S|��L�����οB�<�$=��?�7?�>B>�Ӭ��h�Xл�4��[���'O�>j*�=;{z�O����?6�2��=�7<��C� ��?N���&��>�Pp�(�4�Uvc�P�&�H)b?Qн���.i�?��P?�x��c4�e�0=�<�#�#|�>1V��C3��\��9�&=�y����=��̽>��Z7p��C>p���4����=�սI=��>s�c����;��L       split_indices[$l#L       A                                                                                                                                                                                                                                              L       
split_type[$U#L       A                                                                 L       sum_hessian[$d#L       AC��B�AC�z�A�@&�@B���C�Lp@W9FAӷ�?��B?�X?B�
.@U�A�[5C���@I AÎ�B7�5B&?��?���A05*@��B�jC�r�?��?���@9�KA�^�A�/xA���A�ԈA4��@�7�@�2�@���?���Bg%�A3�`A�'C�+�A@"KA��A�s@p�%A.�/@ţjA���@8�fA+�?̀@�@M6?��@L�3@~�@@��PBP�sA�:@IL�@��?��@[v.C�t�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       65L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       G�7x�;SA���)f<�ڒ�-<�hU�u04����<�Zx=>���F6>��ڽ��]=����ɪj��K�L8 >j
<��o<]�H>����?����>%�����">�>�dm�(�w��8=�7�z>5p2>�#W<��I��Z<�'>)����>�\d�L���ET�=0�!>�Y��#r>����PX�(���;��n�>(��Y>|�'>�a><�T��[h>�H�>Rh�/�>��<<>cr���>�ޟ��	��O��?/Z�=
A���:P>�F=��e��ߞ>9����L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       G                                    L       idi}L       left_children[$l#L       G               	                  ����            ����      !   #   %   '   )   +   -����������������   /   1   3   5   7   9   ;   =   ?����   A   C����   E����������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       G>�;�>���>�Y�>���?�+>e�?	#n?ēf?L�F?;(�?T?    >���>Z�<^��?��z    ?KK?iW;>�	.?&P�?*:�?b>>'�Z=4'�                ?�T�?#�D=�@0?��?�T�?p�}? w�>�T?�^    ?ť�?R�+    ?'�H                                                                                                                L       parents[$l#L       G���                                                           	   	   
   
                                                                                                     !   !   "   "   #   #   $   $   %   %   '   '   (   (   *   *L       right_children[$l#L       G               
                  ����            ����       "   $   &   (   *   ,   .����������������   0   2   4   6   8   :   <   >   @����   B   D����   F����������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       G?�2��8��>�@N��x�?��N�4�@��ax���>��=��=צJ�P7����?U�v�u'?m�8�_c.�:Z>`6�GϬ��-^>w[F�!.��B��=���Ja\�
�X>�ʿ�I>��ڿf6�>�Ӭ�4D�|a��-��<lgA�u��?���?@1�=�����@=�y��zF�I�F������d=>����5=��~>��=bQ���:}=���=|�RS=�<H;dwV��'=�����r�yz>Rl�<%�C��a=>�T=����X=^�P��rL       split_indices[$l#L       G                                                                                                                                                                                                                                                             L       
split_type[$U#L       G                                                                       L       sum_hessian[$d#L       GDND�AcSC��DCny@��A��BJ��C���B���Bp��?�m�@��@,^�@��KBC�C?���A�F�C��;B�OW@�trB9��AZ�@8�4@O
?���?� ?��^@oJ�A�owA��A&��@�L@�+3C�h�AOqBT�@�M�?��A�E�A�n?�ƎAI>?���?ц�?���@�AA�t�A��@51�A�D�@�w�@��@58@��>?���@3oAr�IC��@i0�A�<@	G�BLB�@IJ?꣨AX�@�^�A�#�@�)?�b�A6��L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       71L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       A8����K��=�0e<����r>��ﻯ#:_�>�@=��H���>���<��۾�z>2w��B�>͏x?#=���Ie�>jE�^˯;���>9�>���>}+��� 3>���>kf<�5����p>B�D�n�����?�F=�s}��r=B%h��L�=��>���<��;>�������aN�?n�����=���;�N�>͡@:֕O�g�?�34�>Y�佪K=�����v5>��B>yѾE��G� �>����E�KL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       A                                 L       idi~L       left_children[$l#L       A               	                     ����         ��������      !   #   %   '   )��������   +   -   /   1   3��������������������   5   7   9����   ;������������   =������������   ?����������������������������������������������������������������L       loss_changes[$d#L       A>��F>�(?!?)]_?)��> �T?.y>��5>Ȩ�>�4�>�l�;��     ?8�?�P�>���        >#@;�@>҉�>�B�>��=D�x        ?0��>���>��p?�<>�9�                    >��>�iD?M�&    >�e�            >�F�            >��l                                                                L       parents[$l#L       A���                                                           	   	   
   
                                                                                             $   $   %   %   &   &   (   (   ,   ,   0   0L       right_children[$l#L       A               
                     ����         ��������       "   $   &   (   *��������   ,   .   0   2   4��������������������   6   8   :����   <������������   >������������   @����������������������������������������������������������������L       split_conditions[$d#L       A?� ܾw�>��l?�����g�?�r�>�#���@!�|�'��?z>��;�ʡ�{�*?��{�,�m=��*>^?@1¾���=���?�NV�0�"�,�m=�0�=���fx��~� ���\?���>ׁ�=h�f�6|R����<^>"�!?/��5 >�i���[�>��h=�[�;���=��_@6�@��/0>3Q����?��:ߑt=���: ������W�=�����ZJ��׽��@=�E�=�w�/���ż��=��l�mG'L       split_indices[$l#L       A                                                                                                                                                                                                                                               L       
split_type[$U#L       A                                                                 L       sum_hessian[$d#L       AChH�CK��A�1C��BN�rAL�A�`�Cv@���A,�B#q�@�qs?ȠJA4z�AGCջ?�/�@M>C@T�@&�mA3DA��AD��@B��@nBb?��A�7@�;@�SB�GA�(�?�m?�'�?��?�}%@c�@�4�A��@�)�?�k&A1a?��	?�|�?�o�@�R�?�t@r�b?�&@!�B��o@:[AW��APʔ@�@y�@Ĭ�A��j@@�@)j@��b@�ba@�Um@�A?�"{?��L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       65L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       5:3�����!=ك��a���.(=��>�\<�v���>��q��Xr� �,>"��k8>�v�.�?��i�׾���>l�����>�i�<��@�Ʃ�=�B>L�4���?kcj>Z�.���;�p���9Ľe|��R���k>��'��!���z>����g�?	�P�!��>F>�F�;"�����\=�P�>��<'�"��YB>�3;'��>Ĳ�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       5                           L       idI L       left_children[$l#L       5               	   ����   ����               ����            ����   !   #   %��������������������   '   )   +����   -��������   /����   1   3��������������������������������������������������������L       loss_changes[$d#L       5>�>ܼ>HG>?#��?o._>�@�    ?A9    ?�2R>���>�}�>���>��z    >��f>��4>�G�>h4    =��>x�?r��                    >��?Ifs?
l:    >%9�        >/��    >���>vH                                                        L       parents[$l#L       5���                                               	   	   
   
                                                                                         #   #   %   %   &   &L       right_children[$l#L       5               
   ����   ����               ����             ����   "   $   &��������������������   (   *   ,����   .��������   0����   2   4��������������������������������������������������������L       split_conditions[$d#L       5?ܭ��j���)B>�m2�g�D?��=�n��m���[��?�C��v�}?�i�?B0�>�C�f���@� ����.��=��?,k!�Hn�-8M��eh=Z�=u�?�m6>�;�?m�8?V����Uܽ�q�1��(�N?�L!�{?n�X�)�ڽ��>%i��BE=�T=��g:Cཡ�<=��>!�;IF���(=q:I-o=�	gL       split_indices[$l#L       5                                                                                                                                                                                              L       
split_type[$U#L       5                                                     L       sum_hessian[$d#L       5C��C�@�A�9A/C�/4A���?���@�>�@L>�@ի�C�؅@���A���@]p~?��@�N@�j�C�n|@��)?ɠ�@J��@�%�AE�5@l,?��?�H"?��{?�Ƙ@(q�BBҁC�,?��@;��?�5?�{@��e?�Y�@���@Ғ�?�@(?���B�LA@��@��4C���?���?�6@v�n?��@{?a?��S@�@��L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       53L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       -�)�;:۾";������J�S����9�<K���X�b�=`��;�X�>���=�/��0�����=<z�%�>]��=�X98��>��=�VȾ�lU>�I���޼��⾣1�=�;�;?�>����>Ţľ礰;�]>�td��4�>��z=P���>�<�>�����s>a�<Y�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       -                       L       idI �L       left_children[$l#L       -            ����   	����                        ��������            !����   #����   %   '   )��������   +������������������������������������������������������������L       loss_changes[$d#L       ->w7M>d�>a%�>c�    >a[#    ?�>��D=��>�I2>�r5>�X?>�](        >rp�>_��?{��?�I�    =�w$    =�w�>t7�?{�o        >4�d                                                            L       parents[$l#L       -���                                               	   	   
   
                                                                              L       right_children[$l#L       -            ����   
����                        ��������             "����   $����   &   (   *��������   ,������������������������������������������������������������L       split_conditions[$d#L       -?
�@,�=> ݼ?ܭ���q&��N�ԫ�?�C�>��F?���h3�j���.��;�*�?�i���5�<`>��P>�t�m��i�{>�f=�DW���f?$n�Hn�-8M���A=#־��>���(��=�)��
�j:�o�=�����$>��<3-���K�;��=�����h�=��bmL       split_indices[$l#L       -                                                                                                                                                                  L       
split_type[$U#L       -                                             L       sum_hessian[$d#L       -D~�D;�AP�ADȬ?�/A'�@#��C�?A�#�@h�@ۆ�C���@���@���A�:�@"�d?�Ə@Q�Q@eUA��C�c�?���@,&?�Z@O@۠�AJ��?�,�?�C�@�7?���Ay�@�e�@�)YC�C#?��b?�h�@�Q?�{}@�'2?��@���@�Ou?�Hm?��L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       45L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       M:�5#�92)<ީ��z(�����w]=�$�=�̾��>.�r�A��<eX��s�>�S{<���>B�S�m���L���.<���>ۀ�ѥ�<�&�=y߽����$���>�Uʽ^��>N�&��i�>x2�������>I\>U�n�Qi
=z羾lӾ���<T�>3\�?k9>+�J����>�$'��A�U��>f:X=�>�m�m�¾��>��W�_>�f��;�=�
��JT�=��>�6�>B���Vp��=�r=��N�6�>�����=2�:">>�Cž��F>9�6�G����>�';���L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       M                                       L       idI �L       left_children[$l#L       M               	                              ����������������   ����   !   #   %   '��������   )   +   -   /   1����   3   5   7   9   ;   =   ?   A   C������������   E   G   I   K����������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       M>�w)>� :>�p	>@>�Na>��?��>N�9t� >���>��>�{"<�@>�5�>��                ?��    >�i�>���>���>�)�        >�ƀ>^��>?ψ>�5}>l    ?�>Y/>��.>�pB?K�>��>*tD>�4>���            >��>O?)>�z�=�͊                                                                                                                L       parents[$l#L       M���                                                           	   	   
   
                                                                                       !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   -   -   .   .   /   /   0   0L       right_children[$l#L       M               
                              ����������������    ����   "   $   &   (��������   *   ,   .   0   2����   4   6   8   :   <   >   @   B   D������������   F   H   J   L����������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       M��8��q�1��������Ǿt�>Y�]�?��P���? E>�n�̾�%�>�4`<��|=i�d���Ž�n¼����^p>��@#���۾�?�r$>����0���� =X˶>���?���@-�g�����7����@*A�?����x?��|��m|?��g?���>^�>2E=M�����`=���?�E�?�J�=,�<3wA=����B��eN=�H��[m=�ѽ`j�<���r��<3��=�t�=i�ý��(��<:�<󗑽-6=�.v��|��_\K>
�C��,T=^5;"���=��/:���L       split_indices[$l#L       M                                                                                                                                                                                                                                                                                      L       
split_type[$U#L       M                                                                             L       sum_hessian[$d#L       MCd}�B��,C��@��HB���B���BXK�@"��@��l@��B��B��|@G��AB��B'�Q?�3_?�,@�[?��G@��@�]B�A�*B�h�Az��?ֶ4?���AD@"I@�-�B	��@j�o@D3B�_@0��AYA�~B���A1U@�@bA�o@�؁@J�?� �?�q�@�-@wA��Q@`�@?�ҪA�I�A�|�?��N?ɝ�@��:?���A/�dAg�Bw��@PW�?��6@��\@��?���@�_@M3�@���@��@��@C�0?��?��'A��1@��@�?�:�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       77L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       +9���,u�;z2�~Ԣ={�:��o>�������:�.#��a�>=�����=T��<��¾�o���<<��>5�ݼ�'m�.2�<:��>��d;�Ƚ�z�>���>i�=�g>�־y�H?Ag4����~�8>�S(>(�(m�>���V�0>N&?������>-!����>��#L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       +                      L       idI �L       left_children[$l#L       +               	   ����   ������������      ��������                        !   #   %   '   )����������������������������������������������������������������L       loss_changes[$d#L       +>��><�~>q`>"z�=�>�>P�    >5g8            >��?6i�        ??�?$��?%�?dW?o�?ʝV?/�	?�>�RB>���?�2?I)�                                                                L       parents[$l#L       +���                                                                                                                                L       right_children[$l#L       +               
   ����   ������������      ��������                         "   $   &   (   *����������������������������������������������������������������L       split_conditions[$d#L       +�M��?���@7��?sB����?|�G=��(�M��9�����A�=ckо����j;��ܝ==)��y�7�cH�>=W�����=m�z�\f��X��=�8�¥b?,	�D�=(�h���,>hr�	wǽ��>��=/L��J=3nx��Ʉ=w`�>7D��q=O�ռ�W=���L       split_indices[$l#L       +                                                                                                                                                             L       
split_type[$U#L       +                                           L       sum_hessian[$d#L       +C�YzA�C�H|@��	@
��C�*B@q@��4?�gV?�M?�p|C�<IB���?�_�@F<lB�@C��EA��6B& -B7BQI@�f�C���@�ҨA�*�A�T]A���@���A���?�BJm?���@�<Aك0C�w@3E$@�0A�YA?��Az�@H>�A*V�AAuL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       43L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       9�o�/;6ګ��X�<4���Z�D<f��j�,;���>�/4��c�����>ruG���=�&��j<���jN���?-9��֒�>%���`ܾ�.>�u��nV�1�>v����w�<i>���Y��8�=�>&�?KA ;pm�h�?��<���>�W佗���Ru����<<:B>�v�P��>��>'$7?��׽z�v?���v>-��=F�-?$&O���> ��L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       9                             L       idI �L       left_children[$l#L       9               	                  ����            ����      !   #   %��������   '   )����������������   +   -������������   /   1   3   5   7������������������������������������������������������������������������L       loss_changes[$d#L       9>p�I>u-k>j�w?�$??5>4b�>�.�>�5?���?vn�=Z�    >�wh>&�}<�P�>��t    >���>\@?�?���        >d�<�4                >�
[?Z�            >�^�?i�U?�@>��?]�j                                                                        L       parents[$l#L       9���                                                           	   	   
   
                                                                           "   "   #   #   $   $   %   %   &   &L       right_children[$l#L       9               
                  ����            ����       "   $   &��������   (   *����������������   ,   .������������   0   2   4   6   8������������������������������������������������������������������������L       split_conditions[$d#L       9?�2?|�G��>?z����=�?�H4�4?`�R>l���Ⴞ���=�y�=���P7����@�?�r����U"\�0Zܿ>G�ڢ��j?@1¿y�1�L=��=�9kS��@
pw@Q�?���<(z=HK��7z��0���u�O�6�E�=��߼�U��|�}����;a߃=����z̍=��?=H��>�#i��NG>6@��F�=Pc�<n@�>D�ƾU�=b�L       split_indices[$l#L       9                                                                                                                                                                                                             L       
split_type[$U#L       9                                                         L       sum_hessian[$d#L       9D�7D ��ApWC��B��@�N@��`C�ß@�==BnL�@��1?�S�@�Lh@%��@��C�/�?��!@4�F@k�4B"�A��w?��H@h�=@/�?@B��?��?�Jx?깘@S�QCԸkA�x�?�G�?�\�?�{�@#j6A��_A��@�{�Ab�+?�w�?�|�?��a@<�Cӱ�@a�Ag�T@Lj?�y�?�Z�A���?�ݴA�`f@!-B?��@`��@ =�AB��L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       57L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       G:\�i��
�='k1���þ�n=��R��{ᾧ�::��B��9�=���۴�>	j㾂��<�Ȫ>vE��J&h�/i��<�>�X����=�����q>���=�V���L=�l�n>��滉��<�Hp>��@���0>OfX�S��>;sp���-��UP��l-=��T>����v�����r�=��>��A�Zam=���=��s>�WC�\�<�>0B�, ���Լ�#;�5�>�)S��<=n ����2�\��>j��K����b�=�F��s>4���=�TF>���;�C�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       G                                    L       idI �L       left_children[$l#L       G               	      ����                              !   #����   %   '   )   +   -��������   /   1   3����   5   7   9������������   ;��������   =����������������   ?   A��������   C   E��������������������������������������������������������������������������������L       loss_changes[$d#L       G>k4|>�Ch>^?�>��5>�`>�7�>���    >�Ax>�l,>�}f>���>�X=�K>dQ�>��>�"2>�Dy=��    >Y��>ua<�.0=\<0>��B        <���>�}t>�7    ?_�>m�z>��            <�@�        <�	                 >0s/>�d&        >���>���                                                                                L       parents[$l#L       G���                                                     	   	   
   
                                                                                                                 !   !   %   %   (   (   -   -   .   .   1   1   2   2L       right_children[$l#L       G               
      ����                               "   $����   &   (   *   ,   .��������   0   2   4����   6   8   :������������   <��������   >����������������   @   B��������   D   F��������������������������������������������������������������������������������L       split_conditions[$d#L       G�K�l<�h�>� ۿ���@	���oW2������z�Ծ��D@=ؿ3�r�(ڸ>��X�N���S^>7H0��pv@��=���@P/����$���{�Z2Կ �b������B>6$���i忄��>��2&-�>��=m�=`��F�������Z=��=�>�rk������#�<�l=�(O>cU����<��=�h�?5�F��=S�|�Nj'����7(�:���=�1���|<����	��\�d��t>����<��N��==�����<��U=�h:��L       split_indices[$l#L       G                                                                                                                                                                                                                                                             L       
split_type[$U#L       G                                                                       L       sum_hessian[$d#L       GCa&�C
H|B���B��A�w�B%�!B5�N?��uB��A7s�@��S@ݣ�B
 �@?�4B)��@�[�B�/@���@�a%?���@���@���@a@�ߡA�Is?���?���@ٕB �@T�8@��BӍ�A�@8SF@ �.@��"?�l
@$��?�_?�!4@:�>?�E�?��"?�<
@�О@p�lA�+?� ?��*@�&�B�4?�?��bA 1ZBÇ�@f�@��?�~�?�'�?�A�?�=�?��S?�j(@.��?�YV?�\A�5D@5VT?���?��B'�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       71L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       A�����:m;�w�d`4=o8I;=������f=�Ֆ>^྅�;�Gž����Ώ>�S������K�E��>���>J*��Q����]�<�Iu��<֬��I>��$>������?�=����`����ͼ�e@>�Z���0���8<>�MX<#F+�@�==~;���=������L>�9���ޒҾ�>�xF>��s=o���>(�'����0	�>�˽ݭ��Z��=�����B�U�ܿ7,F<��r��%�>��.L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       A                                 L       idI �L       left_children[$l#L       A               	                                 ������������   !������������   #   %   '��������   )����   +   -����   /   1   3   5   7   9   ;����   =   ?����������������������������������������������������������������������������������������L       loss_changes[$d#L       A>P2?$�>��>��2?)�<?(�n?��]>%Q�>��#>��h>Uײ>���?/��?��@>��= ��            >��8            ?�pt?��o>�$        ? ]�    >熘>ޒ    ?5`>�Z?#�?���>�dH>�>V��    ?9;�>��'                                                                                        L       parents[$l#L       A���                                                           	   	   
   
                                                                           !   !   "   "   #   #   $   $   %   %   &   &   '   '   )   )   *   *L       right_children[$l#L       A               
                                  ������������   "������������   $   &   (��������   *����   ,   .����   0   2   4   6   8   :   <����   >   @����������������������������������������������������������������������������������������L       split_conditions[$d#L       A�ǮO?_�?�p�?�a*?ݙ�?�mO�zz?� ��K�\��@/�P?E4�O<��5j ���8�����mQ=�[?���{���
C;Ծ������f���O�=� �=�bF?+1�>#=��o�?�o�
�H?Ja|?��D?�|F?S�l�=m�>'b�H�<cd�?��(�L�M����=�M���#��K�� u=�)�>^E<�t����=J9c���S>�=�'�һ�%�<�����[��9Q�[λ<�����=��kL       split_indices[$l#L       A                                                                                                                                                                                                                                             L       
split_type[$U#L       A                                                                 L       sum_hessian[$d#L       AC�G	B�C�D�A`	A�#fC�GjA��A2��@4��AvR@��C��@˲�A-�2A�A�~?��?�h�?ݨqAW�?��i@<w�?ַ%C"��CqFA@� ?�W�@Op�@�i�@��@�x�@�Q�@�w@@�7�A�C�|A.��A.ZCff@}+S?�\@�j-@#�?�Sv@Ǥ@=�@�`@0@?�@��&@n6�C�A���@Ҧ�@�	AG�?���C4,kBH�@( ?�$�@Q�{?�Ͻ?��6?�g�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       65L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       -���2<ǰ7��K�<vv�>�X���$���<�ԛ������>����s�>"�<�y�>�H��%޼�"j?4=�>�4�m��ע?8�4=6<�A���)D>m���;�d෺��:>E ��W?����<�DY>�q��S��>���=�� ��}>�P¼3��=3���+\=�iy��SL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       -                       L       idI �L       left_children[$l#L       -               	����         ����            ����������������         ����      !   #��������   %   '����   )����   +������������������������������������������������L       loss_changes[$d#L       ->�f�?9��?8).>�Ҡ>�d    >иI>���>�H    ?�4?� �?e�>��                >?�)?qF    ?�3_?>�O?�3        ?Q�?�    >�4    ?�m                                                L       parents[$l#L       -���                                                     
   
                                                                                L       right_children[$l#L       -               
����         ����            ����������������         ����       "   $��������   &   (����   *����   ,������������������������������������������������L       split_conditions[$d#L       -�.p��X��V@B�9���,�&�?�ͨ@@Vʿ%}�:�.>w[F?EU	?�	L?�|F>;Ž��>��)L>X$�)���f��(�>]��߾�?�!�{�=���EW������i�=lxg�q
�>8z
=D�;��=����~]x=��<��Z���E=�-��W��<)�M8<�K^��	�L       split_indices[$l#L       -                                                                                                                                                                     L       
split_type[$U#L       -                                             L       sum_hessian[$d#L       -DJWCvnC�T�Cpro@���?��aC�]uCl�Z@e�J?�ޢ@��(C��JAU%nCk��?���?�l?�w(@�@ �>C|��A)ڠ?��jA@l CWVA�,?���?�ϚA"8CCr�f?���A%?�ZA#��CS�@y[�A���@��@}Z@��X@�{,Cj��?�ώA�3@�9y@VL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       45L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       :"�>T��h�D=Ȥ>������;����c�,�O>����&މ>ڤy>/>��gL;"����>�y�>&;�
�&>�ћ�MW2�*�w;!e8L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L                   L       idI �L       left_children[$l#L                ��������      	��������      ����   ����   ��������      ����������������L       loss_changes[$d#L       >m��<Z ?Y�        >̰>��S        <	��>�?e    >u�T    >���        >��>��6                L       parents[$l#L       ���                                   	   	   
   
                        L       right_children[$l#L                ��������      
��������      ����   ����   ��������      ����������������L       split_conditions[$d#L       �p��<ߠ(�o�|<���=���;�l�m帾�
�O�_��Ȱ�l��>/|�+'P�
ȿ��Z��i=��>�z�f�K=��T�vh��L�\:A��L       split_indices[$l#L                                                                                            L       
split_type[$U#L                              L       sum_hessian[$d#L       C]�@,MxC[BI?щ?��@�n}CV��@C�d?�o,@�<ECR��?��@8�?�܊CQE:?���?�rA?BCEQ@�ck@� �A=�|C9ubL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       23L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       ��>�M�>{9�b�|�� �[ >{�ӽёr�ð�:}��n7�=��>�w��>�?A>#���#����>{���K];��H��)>�{���d�$/"L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L                    L       idI �L       left_children[$l#L             ����         	   ��������         ����   ����      ��������������������������������L       loss_changes[$d#L       >OE�>�k    >��<H��>�%+=U8        ?0T??:=�	�    >���    =��<��                                L       parents[$l#L       ���                                         	   	   
   
                        L       right_children[$l#L             ����         
   ��������         ����   ����      ��������������������������������L       split_conditions[$d#L       @X�@Gh^=��_@,�=@W�l@
�?j�ܼ�{V���b@
ڬ�Xň���~=�<)��n=�?
X>��l����=����-8:�~W�8�=�-�"�߽E]L       split_indices[$l#L                                                                                               L       
split_type[$U#L                                L       sum_hessian[$d#L       C�fC�c�@�C�@�@~<C�@��+?�ٍ?�"�C�z)@��7@_��?Ò�C�S�@M�@ |�@���?���?��A߸C�X?�v�?��O@)`�?�!�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       25L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       +9��;o����Q��;���;y�2�b�<������2>��r:���>`�ӽ��(=�N��lL<��'d2>�� =2,���;��5=�Bi�v� �>V�������w�>�P�=�Ŝ��7���/P>�$:%^�>��e��V���ד��W+���0>,�H�>�����ߔ;��]L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       +                      L       idI �L       left_children[$l#L       +               	         ����      ����         ��������   ����         !   #������������������������   %����   '   )����������������������������������������L       loss_changes[$d#L       +>]�>M`�>E��=.��?*�>�>���=�    =��H?/�    >s��=�D*<od�        =`��    >$s?<�>=Tx                        >�3V    ?��?I�J                                        L       parents[$l#L       +���                                                     	   	   
   
                                                                    L       right_children[$l#L       +               
         ����      ����         ��������   ����          "   $������������������������   &����   (   *����������������������������������������L       split_conditions[$d#L       +?�2�p����><ߠ(�o�|?�H4�4��z��أ;�l�m�=��=���P7����<j�Hޣ?�Z�<U�i�nl�j��>w[F@
rн�Y=���1�վ�z>�<Ć��V�r��ʿ|���it5=�������i��h���i�=3�����>R��L:�o�L       split_indices[$l#L       +                                                                                                                                                              L       
split_type[$U#L       +                                           L       sum_hessian[$d#L       +D�5C��RAc��@dW�C�ڢ@���@�F;@ �?��@�j�C���?���@�Qw@iM@���?�ǩ?��~@��q?҉�@�f�C�\@.JU@8X�?�7�?���?�t7@=�@^�o?��@r�B@*w@��C���?��?��?���?�#I@(�?�<�@-�@�O�@���C�)L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       43L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       3:G;=+\���y<κ�>��#�@����ذ:���>E������<�����;� <pR���FD>�<ݽ���������b>3@s��7Z<V$S����<oUe��=����ꇾ>>�bc����>z���#>C��۰�>�6=��񖽎v;��&>p���n��a��<���>�tx����<�,v>��4>�L��i�=��>�F�:= L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       3                          L       idI �L       left_children[$l#L       3            ����   	                        ����         ����   !��������   #   %   '   )   +����   -��������������������������������   /   1������������������������������������������������L       loss_changes[$d#L       3>e�?
��>վF>��     >�\>�U>�\�>��=�[�>��>cN>��t>�    >ƸV>i|�>f��    =�gr        =���>m�\= Ҡ>�(y>�^    =���                                >j7�>�                                                L       parents[$l#L       3���                                                     	   	   
   
                                                                                 %   %   &   &L       right_children[$l#L       3            ����   
                        ����          ����   "��������   $   &   (   *   ,����   .��������������������������������   0   2������������������������������������������������L       split_conditions[$d#L       3�1㠿4�J����?��>,�?�ʿ*�V? �}����v�?@1½��@9�0�A0��]\�g�������v��.8��u�;�|2��'@�l?�>���=:�(?�A����O=J���R�=j�7�А=��}�]��������@*5��9��q�;��=�Ľ��z;�(>�=.�\��Kl<'x=�!߼_|gL       split_indices[$l#L       3                                                                                                                                                                                         L       
split_type[$U#L       3                                                   L       sum_hessian[$d#L       3C\M�B��C
A�B��@5�AN��B���B�C�AۣA9@��/@��B�@B�?�"�@�+�@6@�*@ @`�?�|?�/�@G��B�;�@ ��B��@�6Z?�3�@���?��??��-?�@�?��?��"@��@��?�ٶB���@g�j?�:~?�ޜB{�1@�@Z�?��s@f�?��{B�zB��r@��?�+!L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       51L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       G��ڭ�S4=?��҂E��Ea>s�f�0�:�z>��ν>W�;���>f3���r<���1�뺄��=���?t�����B|��Bp=�L�>�qr<N����L[��>3?��^�yٗ=�!�:��<�Ӎ���0 >+��ږ>#0>G�ݾFu�=F	`?��(�v>K��>Q�g��'�=Y�a�xUT��0�>0N/�%�>�������>��#��_h>�2��j<��*?$K�>x������>��>�&��=M��>�W��C=�B�>��I��pO�܏T>��6L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       G                                    L       idI �L       left_children[$l#L       G               	               ����                  ��������   !����   #   %   '   )��������   +   -   /   1   3��������������������   5   7����   9   ;   =   ?   A   C   E������������������������������������������������������������������������������������������������L       loss_changes[$d#L       G>U�?��?q�?5_>Њt?�3?G/�?��=��?4j    ?B�	?�}�>���?(��>��>���        >�s�    ?)��>���>M��>�cu        ?�%?�(>�.=���?'                    ?f!�>X�    >��?ͳ? ��?V��?7�?�n�@..                                                                                                L       parents[$l#L       G���                                                           	   	                                                                                                   %   %   &   &   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .L       right_children[$l#L       G               
               ����                   ��������   "����   $   &   (   *��������   ,   .   0   2   4��������������������   6   8����   :   <   >   @   B   D   F������������������������������������������������������������������������������������������������L       split_conditions[$d#L       G?0\�?#�@?�d�?П���<�2L?�����<�����l�=5���V6>�+�"f;�[>?�V�?nf<���>!Y,�Z��ia�����&� �bֆ�#�����6F�?^�?~ �?���>AA�?^���3���4=Mؽ�;N=C�6�,�j�>JG<m�ڿ)T�?|a�?\Kb?:0?za�?�ͨ?*�4��:j=S��F�=�,Ժ�\�=�Cļ���>g����;�0�>E'g=�3����= F=�Ƚ#ݶ<v�>
r5��=��=ŷ%�ӹ��V =���L       split_indices[$l#L       G                                                                                                                                                                                                                                                               L       
split_type[$U#L       G                                                                       L       sum_hessian[$d#L       GC�մC��B��[C�d6@�9�B&�B�kC���@6�6@���?�pA��'A�3@A��B�]�A�o�C���?�bc?�"	@U��?���@Z�kAz�3As�AP�N?�� ?��QA�B=��Akj�@��C���?���?�D?���@�X?��'AC[@\s_?��QA��@��@���A�
k@ҪrA���A���AQ�?�� @?�?���C��@�I�@�<@��z?�+�@
]l@��>@Iqc@u F@;-@|C.@X�A`�@���@$wg@�n�A��A��Ac�@��L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       71L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       9�g�V;~��)�<W��7յ�B����b;ߛ)>�Q�>-����>^�[�=v�<+����-�>��<��ؾ��>���]�ؼDɻ?x6��ܮ>�N��}ӟ��G8> \h=����Un?�">4�=WԂ�?&>�=��$`+� $3��v>�fh�)�>�!T����;��X��oa>pH���)ʾDee��ռL�<?	^A>6�"����<t<����<A.�|#�"1>Z<�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       9                             L       idI �L       left_children[$l#L       9               	   ����                           ����      !   #   %������������   '   )   +����   -����������������   /   1   3��������   5����   7����������������������������������������������������������������L       loss_changes[$d#L       9>O;�>g��>~��?l��?a�?>�V�    >��3>P?_�c?.b�=���>qb$>�W�>�C<Y��    >�Kl?/��?A� ?;/            >��>�$?AC    ;�%�                >��>���?<&        >à�    >u M                                                                L       parents[$l#L       9���                                                     	   	   
   
                                                                                 !   !   "   "   #   #   &   &   (   (L       right_children[$l#L       9               
   ����                           ����       "   $   &������������   (   *   ,����   .����������������   0   2   4��������   6����   8����������������������������������������������������������������L       split_conditions[$d#L       9>]R>&kh>���>�0��#��A��
v=�B<?�@^>���?{S�x��3S�)!z��={�;�Gо�@?�>��?RԺe�u��<=�^r�X����?��Q<��ݾȠ>Ґ=X�<���(KȿU%>͙�c[:�(�>p�=o�d=���>;�,:�������=�+Ǽ���k��8���u��>$ׂ=[)���;��Ƚ���;g�k��H½B�H=��&L       split_indices[$l#L       9                                                                                                                                                                                                                L       
split_type[$U#L       9                                                         L       sum_hessian[$d#L       9D_�C���A���C�B��_A�L@S~C��t@��0AiVDB���@�U7AH�C˳@���@��?�%�@��AE�ZA���B�@?�zb@um=?�"�A8I2C��B�`?հ�@$T�@TU?�а?�??� 1@�}@�_�A���@�`}?� �B^9@+"A~jC���@��A��DAA��?�b?�G�?���@���@[��?�̓AF;�A��A��N@���A�?�3:L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       57L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       K�5���1�^<��񾃨Ҽ�����R=+��{W��̇> "@�`��<?�2���>��<�I>��.��R����<,G4>�c��&����>����/��=~>�?��=ٮ����>�mE�J��;�1�>%���F�b�e>Y����"=Q��>��޻�2�>�9����=�D�>8{s<I���V�>�׃��:[���>pRC��Nؾ*� >s��UC�uO>�¼������E���D>������'�k>��K>n∿ �?uP>���<��@ �>R��� ��=y�[>� ��4�r=�}�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       K                                      L       idI �L       left_children[$l#L       K               	      ��������         ����                     !   #   %   '   )   +����   -��������   /   1   3   5����   7   9   ;����   =   ?   A   C   E   G   I������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       K>e�>�P�>s�=���>ǎ�?.iB>��        >�S?>u�E>��    ?% />wP�>u�>�8]>�43>���>�F�>�=`?�?�>��>���    >R_�        >���>؝�>�*�>��`    >ɗj=m>�    ?	��?DF�=UV�>�0>�h>�0>��)                                                                                                                        L       parents[$l#L       K���                                               	   	   
   
                                                                                                                 "   "   #   #   $   $   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,L       right_children[$l#L       K               
      ��������         ����                      "   $   &   (   *   ,����   .��������   0   2   4   6����   8   :   <����   >   @   B   D   F   H   J������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       K��8�w��9�e>Ɍ}���ǿH�!�CX<�Ҕ��(��4��>�|�=m���{�b�c>�<�f���>���ݞ��o�>>��6�+����?��?=�J> l�:��*���=�� ����?}��H���&���棿z�d��?� >�]>&An�P��U����>��P?�1?�9���h=�5Ѽ�ߡ��]=�1\���7�M&'=�+�ٙ����=������U�=�wӼ U��IN=���=�T��e�>4��=�V9<:��f��=|���sr<��j>��X�V<���L       split_indices[$l#L       K                                                                                                                                                                                                                                                                                 L       
split_type[$U#L       K                                                                           L       sum_hessian[$d#L       KCY��B��C�o@��@B��A�UHB��@D�?�Z�A�Bl-A��X@c�A�oB�L�@�+�@;VB��A��AKA2�dA���Ab/1B,��B)��?W@���?�/�?��A�HAn�A�A��?�3&A��@s��@��?�-�ApA�@���Ae<B��A(<�A= A�Y-@E�
?���A2�o@�%d@���A' �?���A if@��A��J@��5@x�.@,�L?���?�D.@���AE_@,�p@Y�0?�?G?��^@��Ad��A���@�x�@8�A{�@:��@�N�A��{L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       75L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       :TJ#��;���T�>'+>�e:��f���ؼ��Y>֝��!�:��	�;|dо� ��O�->���>��B:�/ھ�d=�8Žڦ�;�ֵ�T ����6>����P�>>ꣲ;"��L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L                      L       idI �L       left_children[$l#L                      	����         ������������   ��������   ��������      ����      ������������������������L       loss_changes[$d#L       >[��>��
?NB>��>��    >�,�<���>���            >��        >,�m        >Xl�=��    ?X�4?.&p                        L       parents[$l#L       ���                                                                                      L       right_children[$l#L                      
����         ������������   ��������   ��������      ����      ������������������������L       split_conditions[$d#L       �Yt�<�UE�X �>�Ӭ>�b�>	y�Rd���6��Wy> ��Bཫ�/�J�T�,\ ���t>&�Y=�l2=���#��DL~=�w�;n�!���~g��=�2Žz>Ȟ:CL       split_indices[$l#L                                                                                                                L       
split_type[$U#L                                    L       sum_hessian[$d#L       C�A=�JCܴ�A�@�k?��MC���@�&@��W?���?�S�@~�C���?��`@@��@`�??�n�@�Cٝ�@K}?���A�GxC�y?�^3?�8�@z�A^�?@;C�R�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       29L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       ��q�:4����;�ξ�P9��>��T;� ��H�>��Z=��l��kE;���Z]d��;=� [��ޙ=�F9���O܆=��lL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L                  L       idI �L       left_children[$l#L             ����   ����      	      ��������         ����������������������������L       loss_changes[$d#L       >G�s>9U�    >��@    >��[<�
�>D:$>jʨ        ?��>��/>s:k                            L       parents[$l#L       ���                                                              L       right_children[$l#L             ����   ����      
      ��������         ����������������������������L       split_conditions[$d#L       @,�=?�4�����?�*F���?p]�?Nv��K�>���=�.m<��O�dF4�`��?OB��{<՚����=0�8�U�yo<޴�L       split_indices[$l#L                                                                                     L       
split_type[$U#L                            L       sum_hessian[$d#L       C��C� �?��C�_�?�O C�S#@>�C��oA9�?���?��AI�xC�=A��@[�@��p@̔�A�m�C�-@�p^@��L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       21L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       M:�;=Q��[�: �>vv���X=#�b<��N��D�>֘�=����!��&�D=�R��"�;�s�>�EоĶL�S�S��>����־�/�=Î���X�>�=_���F>\�Z= �%��>�ڗ<�e��$�ž�vľ��>��8=�<��E�=�}�>� ��{>l޾�>���:��	�#,>�P���E_��nK=��>���;�+ϼ���>ՐH�s�>��>Z�3����*�B���y��{��]��>�W�<��ھ S�=�V��i�=��ؽ~��>~��=�"�����>?���!�վ-�>;�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       M                                       L       idI �L       left_children[$l#L       M               	            ����                        !   #   %   '   )����   +   -����   /   1   3   5   7��������������������������������   9����   ;����   =   ?   A   C����   E   G   I����   K������������������������������������������������������������������������������������������������L       loss_changes[$d#L       M>`��>��o>�t.?�h>��->غ>�>��a>i�    >��>6t>a��>�G�>�TQ>{�)>*�(<���>�O>hf�>ix>�x�    >�>��h    >��i>���>:��?�Pf>�3                                >��    =��h    =��j>w��>ս�>���    >���>{1p>,`�    >�                                                                                                L       parents[$l#L       M���                                                           
   
                                                                                                               '   '   )   )   +   +   ,   ,   -   -   .   .   0   0   1   1   2   2   4   4L       right_children[$l#L       M               
            ����                         "   $   &   (   *����   ,   .����   0   2   4   6   8��������������������������������   :����   <����   >   @   B   D����   F   H   J����   L������������������������������������������������������������������������������������������������L       split_conditions[$d#L       M�d��|�j?\Kb����h�$�I�">+��?[/D�� g> ��L�~��5l��v����?���P}��?ƃ��UQ�!�G����*˾�J���v��j׳=��#����>uZ=�kv����<�=�l�<<��Ev�������=�D=�ؽه���P=����V=���"���(��GX?���=��>���>�q�?v�=��@aܻ��> #_��+=-o=�M�J@�L�P���+���º��O>�#;��ӽ�<<�g뽋��<�U����=�ؾ<�\��ѭ�=fcg�Bg�O��=`�9L       split_indices[$l#L       M                                                                                                                                                                                                                                                                                        L       
split_type[$U#L       M                                                                             L       sum_hessian[$d#L       MCV!�Bɤ�B➄B��A�7B�R�B*�lB�6U@ʳ�@e�A�?zA��Bxh A�QAq��BG�@�'�@��@@?�tA�DK@�5�@lA�(BS��@U�?A��NA6e�@mVXBW~A!�@?:�?�*�@ Ӧ@t�?�6b?��?�|�?�6!A�MR?�o�@�|?��@rl�@�A���A��L@EA��@��@���?���@�BA/�@���@��@.%�AhfA2??�w�@J=)?���@@1�W@&T�AX�A�a!A���@�e�A�G�@V_�?�3b@�G"@OH�?�Nf?��K?�UxL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       77L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       -:^j����=����%��8(#@�So�> Tq��k�=Y�>��ɻ�q>�
K�,�;>��"=��o����f3��	9>�a@?E�V�����ݎI��
���=���<c�>����i�ھj>���=�P>�v��fH���	=9��>t,���f�x��>����җ�?ꀾ��6:96��>��L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       -                       L       idI �L       left_children[$l#L       -               	                  ����   ����   ��������      ������������      !   #   %��������������������   '   )����������������   +����������������������������L       loss_changes[$d#L       ->Z >�Z�>m�;?�?���>���>��>N�h?T'�?0��?F>    >fa�    >��        =@yP=�P`            ?T:>TI�>ө>�u�                    ?���?>                >��2                            L       parents[$l#L       -���                                                           	   	   
   
                                                                 %   %L       right_children[$l#L       -               
                  ����   ����   ��������      ������������       "   $   &��������������������   (   *����������������   ,����������������������������L       split_conditions[$d#L       -?ܭ��g��T�z>��P�a�b�h88�*��?��?T�?P#��jX<=�Z�9ND=�"�;�A:������?�@^>�A�>m5��vȾ���g�D>�Cu�%bF?��P=�e�2���h>.�<�v`�[���b���'?<^�/=��ڽ�����=�둽��2>�4����9^A����=-��L       split_indices[$l#L       -                                                                                                                                                                   L       
split_type[$U#L       -                                             L       sum_hessian[$d#L       -C��MC�9�A�|�A'��C��~@瞠A)�@�z@�d�@G>ZC�m?��F@�l@85AW��@g��?��@'��@F��?�k?��I@��C�=�@j��@KA6a}@�;?�c]?ʄy?�?���@���Cˏx@"�?���?��?�k|AP�?Їi?�k6@���A	#�C�FX@�� @�� L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       45L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       A�|} ;�Ѥ�q��;5
:>�nO=����C��<x���	>�K��"v<�v�Ӎ �$H=Њ���޾��(���>�9�J~D>;q����*>��(�NZL��o�3�q���?��<��P<�Ⱦ���;��쾵�y?�=W�>"-��A�>�k��%�J�i
�>+��?v�=����'�F>�uݻ���E��W��=5%�=�O��8������ʾ�"s>^Q�FS>�n=ʱG���.��[d��7e�l�->�3��J�>s��L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       A                                 L       idI �L       left_children[$l#L       A            ����   	                                 ����   !   #   %   '   )��������   +   -����   /   1��������   3������������   5   7   9   ;   =����   ?����������������������������������������������������������������������������������������L       loss_changes[$d#L       A>8]>��=?Z�>Y��    ?0��?���>à�?M��>�Z�?5o? ��>V��?C�p?/�t?O�>Ac    >��>�5@?&�<>�N->��        ?���?���    >�W>�/q        =�            ?by>l��>$K�>`tn=�g3    =�u}                                                                                        L       parents[$l#L       A���                                                     	   	   
   
                                                                                                     $   $   %   %   &   &   '   '   (   (   *   *L       right_children[$l#L       A            ����   
                                  ����   "   $   &   (   *��������   ,   .����   0   2��������   4������������   6   8   :   <   >����   @����������������������������������������������������������������������������������������L       split_conditions[$d#L       A>�,�>��ܾ�>��*=��Ƽ��$>xn��(�>��=�{�?O���<B���@���C���?�ٳ�#����2?�o�H}E�g�$?�6$?=��w���4C���>��>5��X���29D�ؿ�;/�>5q�>�B<���=B�j�_������?:rT�4��Z�>"���
���Ik!>��	X��m5ݼ�n�<Y`f=���"DV��ʽ;���揾=�d^����>u�<�;#���8����u���O=��f���=�A(L       split_indices[$l#L       A                                                                                                                                                                                                                                         L       
split_type[$U#L       A                                                                 L       sum_hessian[$d#L       AC��C�U�B=��C�V�?���A��4A��[C�/�B��@Ǚ�A���AB��A2U�B�	0C}[ B�b�A��?�Y�@��A"�@���A��@pU=?Ֆ(A�B��@���?�ŴC|)�B�#l@g�]?�6�@��'@u/?��*?��A\@��@7K�@�Ӊ@�??�5@/:�B��2@r��@��@!��B�CW��A�7�B��x@�Q@b�B@�]�?�C�?�k�@f !?��?�ھ@5�@b�"?�n?��?��*?��HL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       65L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       5;�<e�U����;��x>I��xaD��h�<��e��a+�K+=>��=ȇd��e���'�=1<�;�� >b�$�Q?k>���>��¼�����#ܽ�Cվ ��=��$<|�4��㉽��f>����Df;��ƭ>���;�=���>�Pu���'=2 �>Z9��v��0=� �=�K>��H.�>.���������>K��Q�>�ڢ�C�6��,s=��L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       5                           L       idI �L       left_children[$l#L       5               	            ����   ����   ����                  !������������   #   %   '��������   )   +   -��������������������   /   1   3��������������������������������������������������������L       loss_changes[$d#L       5>[2�>�I^>p8�>_��>�w>���>�=z>�<? {�    >p��    =��    >Oǭ?L�>�N!>��=��=�CH            >��>��2>~��        >�>��=�BX                    =aw>��>��c                                                        L       parents[$l#L       5���                                                           
   
                                                                                 $   $   %   %   &   &L       right_children[$l#L       5               
            ����   ����   ����                   "������������   $   &   (��������   *   ,   .��������������������   0   2   4��������������������������������������������������������L       split_conditions[$d#L       5>��^=��Z?;��S����o�5j �:M�?�d��s�}>�@<�y?���JA�_]� ǰ=�6�@ �'?�.�̡���^<�̈́�?s��>���>s4����G���%?�aO=�7:>��;m<�g>����=�?ƄT?v�?2R�;��<�=Ɯ>ow�p8\=Q�þ�$��w==9&Ѽ�.�=��)�k!u��h�=��L       split_indices[$l#L       5                                                                                                                                                                                           L       
split_type[$U#L       5                                                     L       sum_hessian[$d#L       5CR~]C:�A�}�C2�@� @�]�A��:C%A]�i?��Y@��J?�c�@�E@3�A}
�C�@��A:|I@8�@��?���@[u<?�)�@�A9��C��@K��?�~B@��S@�n]@��4?���?��Y?��.@@7?��4@W�@��]@zD�B�n�B+�T@D��@$��@u��@�@n�?��?��?�:@��2?�D�?��@P�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       53L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       3�÷���=�;h��H��<�@��K�<!`.<�I1��b�%5Y=���=Qr����?60�;�Ѿ&�>zg���I����>Y�����Ǽ�[�?����5<�6��Ih<�߾=K�Q������¼�&->5p�o�����2[>T	<k�i�` �>B�پ�S¿2����e>�ҝ�EK=����:��%#=(��?t7:,�C>v�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       3                          L       idI �L       left_children[$l#L       3               	            ����         ����   ������������������������   ����         !   #   %����   '����   )����   +   -   /   1��������������������������������������������������������L       loss_changes[$d#L       3>G�8>#��>bq�>B�x=�2?IYz?��4=�.q=�    =��>?L��>��
    >�                        ?�    >�n�>e�?�>���?+T=    >%��    >���    ?M�>��?���? b                                                        L       parents[$l#L       3���                                                           
   
                                                                     !   !   "   "   #   #   $   $L       right_children[$l#L       3               
            ����         ����   ������������������������   ����          "   $   &����   (����   *����   ,   .   0   2��������������������������������������������������������L       split_conditions[$d#L       3��8\?��Ozo��l&>�ŵ�[��M��>�� >M l�F@=�u{�]|?n��>Z�%?��ֽ ��=/���X��<�=�����i��]�H>2�<?�{�J��?~(P?�i�=�k�c?d���-пU�t����>k�n�?�j@^e��f�=i�������Vg��5�>���)�<��G��V����<J��> %9OTQ=� :L       split_indices[$l#L       3                                                                                                                                                                                      L       
split_type[$U#L       3                                                   L       sum_hessian[$d#L       3C�|DAEW�C�Q�@�M�@�bCA��C���@/=�@���?��&@L�tA���A>�	?晤C�	\?���?��`@]�Z?�)�@�?��A��a?���A	�@k��C<5lCU�LAz�_?ף@�_2?��@$�?�;HC5�|@�~A�C9LJ@��A'�@��?�h�?���?�79B�c�B��M@��[?ǒ�A�`�@���C/�A#�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       51L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       +�k�;;=���\N> ��9�I=�%>;�ë�g�>�ɚ��������C�Z>�cᾆ�E;)
>��=�>�ő��ؚ?O���]>@�t�cI5��>J���4 �< 	G�K3=t�.��d˾�2<�+yu>ŗ���=<;쾣�Q;��~>�bؼ��[��Q��˪Z��L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       +                      L       idI �L       left_children[$l#L       +               	                        ��������   ��������   ��������      !������������   #   %   '����   )������������������������������������������������L       loss_changes[$d#L       +>0�p>2E�>N[i?�k?(>!=���>���?&�>d�>�A>�	�=��$>G��        >81        >r($        =�:�>6�            >u`>��>�=    =c��                                                L       parents[$l#L       +���                                                           	   	   
   
                                                            L       right_children[$l#L       +               
                        ��������   ��������   ��������       "������������   $   &   (����   *������������������������������������������������L       split_conditions[$d#L       +?
�@5��>���@�@@�n>r�,>���@
�1�	l�'��@Q�?�9����>o!����?|�G>
<��#�O�+��jS>9,ǾތF@SR���_ ��|!=s*Ͼ6��?z����=�<���>��P����M��=�F�*��<aႽ�;�:�1=�����Խ��t��f��JL       split_indices[$l#L       +                                                                                                                                                              L       
split_type[$U#L       +                                           L       sum_hessian[$d#L       +C���C�T�A2� C�H"A!��A!�@v>C���A,��@u�@�<�@�R�@���?��v?�C�/[?��-?�j�AY8?��@a�@`��@/��?�hn@E�	?�x@8$�C͘?Bd��?���@��@
�s?���?��a?ֶR?���?�P<C�k�@�#|BP�E@���@��2@��L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       43L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       W:i��=	`��*;<1�.>����5�=;긼Ϊ=��X<F��>�J���=��>Ƞ��J�/;�����>�FE=o`,��>��>��> � �b�ؽe���*�>|N=��>������=�|μ�F�>�"�� �����=�
c�t��=[�>���;�T��J�=��c�$W|<��!=�����<����O>� r>T.��y�>I�%�~0�;��#�s��7Y�>�J��5�׾��>�s>�&߾� )>3�1;�켼)��bUJ>�G�@W�>
S���9�mW>eoý6�=�ʾ],>)U�� �Z>*`F��BJ>�8�"�w��!̾�׃>� ��O��L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       W                                            L       idI �L       left_children[$l#L       W               	                                    !����   #   %   '��������   )   +   -   /��������   1   3   5   7   9   ;   =   ?   A   C����   E   G   I   K   M   O������������   Q   S   U��������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       W>P(�>w]�>���>�l�>��>�^2?�f>�c>���>}��:پ >�-�>w�>$l>��]>�in>;�d    >Y$p>1�>IF        >�)(>�� >�B�>�
{        ?~��>��>�վ>E�~<y��>���>�	e>Y'=N��>�c    >�M?/�=c?>�K�?��>f�4            >���>M�>�8K                                                                                                                                            L       parents[$l#L       W���                                                           	   	   
   
                                                                                                           !   !   "   "   #   #   $   $   %   %   &   &   (   (   )   )   *   *   +   +   ,   ,   -   -   1   1   2   2   3   3L       right_children[$l#L       W               
                                     "����   $   &   (��������   *   ,   .   0��������   2   4   6   8   :   <   >   @   B   D����   F   H   J   L   N   P������������   R   T   V��������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       W�d��d�?�9:�zH�?��?���?�&����<���>��6�ABؾJA>�#�>�$�?��?[/D�� g=�TS�J���=^��|a�=���=@��@UT�Ei�>h����`<#>�?K9r>�����߿0�뽢Q�����T�?r��>�8�����=�כ�e�n?�(@-d����>� �>C�l��=�^c>
 E�n5@�l�m@O-����:��*����\3=���Yޜ�����q�=��!=�����e=.��+�]����˅����=����f��=&2d���9P=��u�"A�<�I����=K3��Vl=Ls����=Ԫ��C*���[½�5�=ɚM�y�7L       split_indices[$l#L       W                                                                                                                                                                                                                                                                                                                           L       
split_type[$U#L       W                                                                                       L       sum_hessian[$d#L       WCP_jB��Bڵ�B�7cA�F=B�<B�Bl�A��A.��@�U0Bf@A�o�@ddB �DBS5a@ʝ4?�R	A��^@��@��@b?�P�A�#�B$.RA3��@�@�?�$
@�_A�/�ARnBC�	@wex@���@��@Q�OA���@J0�@�@ �S@d��Ag;/@/�A�czA��*A!�G?�"�?��@>�A>�A JA0��@�eB3 Y@���?��5@1�^@��?�(?�@p?��I?�9@��A�N@�/@3�?��9?�V�?���?��@�%@���@�ɷ?���?���@L�nA]�AA��A>i@ظ2@T��@ym@�� @�m@�h^@���@�`L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       87L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       O9��ܼW�=�G�ܙ�� a=�:;���&��2$;����S�>/e���=��G�B �=���>�|M9*�����=��? �l>xA>`���y>�$��"y���f�K%��fU>p�M����=����M�:������>���?�
>���͊�>w[}��H>��	=Q:��E�>ӕ�45��SK=dh7��BL>��!>z �~�=�@�������>�ӓ�4�P�'�>D+��k?>(�A���n>���o>(~׾�v2?"-�=��/���:>��$�*+ʽ�_�>��=���^��k�>���$��>�	��"`>^�WL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       O                                        L       idI �L       left_children[$l#L       O            ����   	                           ����         !   #   %   '   )   +   -   /   1   3   5   7   9������������������������   ;   =   ?   A   C   E   G   I   K   M��������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       O>f�?Yd>Ԕ>>�     >춚?2b?,#>ǖr>���>�p?�Z?q&=?#�8?'�z    >�Ϳ>Tr >^b�=|o ?P��?/��?���>��?z]�?��U>���>K��>�ܚ?z�?CϾ                        ?:?7�">���>H�@?�0�?�>w �>�q1?���? �                                                                                                                                L       parents[$l#L       O���                                                     	   	   
   
                                                                                                                     %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .L       right_children[$l#L       O            ����   
                           ����          "   $   &   (   *   ,   .   0   2   4   6   8   :������������������������   <   >   @   B   D   F   H   J   L   N��������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       O?0\�?.�?�d�<�h��F��ǮO�L��?�\>D�?Ja|?9��9O�AE�j{��*�=��]>��w�f^?[�,=�k�6��HC¾V6� ��;n�?O>>z.��D����>~�?�f@� ��:�2�4œ=��5>>?@=*e�[;�?n�>�n�?
X?%�?�g�?t�2?�׿�X>�9־��=��=���21�<�<�ѻ��)�>K��X�a�Iqf=kg��9M=J����p�=�
l�;�m=J1Ͻ��<>B�M<�"���#=�žL4����J>�X��ؽ���=�I��E�Z=�$��=��hL       split_indices[$l#L       O                                                                                                                                                                                                                                                                                         L       
split_type[$U#L       O                                                                               L       sum_hessian[$d#L       OC�G�C�kIB�qzC���?��B�B� �BE�C�@�%A�b
Aט-BF55A�$�A@�?�d�C��@�,@ST@��A�d�A=�nAqQ�Ab|B\�A9��Av��@m<�A~�Cc;�Bc5s@h�?��?���@m5?�QR?���A�NA�|�A	i�@Q��@���Ar�@���@�X@��B
�A!?�	@YgyA@X�?�^E@'��@�:5@�éCa��?��AA��?A�@���@���A���@N�@��*@RIh?�:�?�is?�(�@og~@�i�?���@�v?���?���?���@p�.?��A��@A7ψL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       79L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       #�Y�_��>'/:�0��L�>����yv^�b�>·F��@���U8;���?#����>=��:Q6���ǽ3
<��h>��+�R��f��8����>�jĻ �>�"��d_=���;����+�i�t>����%�;��lL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       #                  L       idI �L       left_children[$l#L       #               	         ����      ��������         ����������������   ����������������         !����������������������������L       loss_changes[$d#L       #>6�U>�v�>��@>�	�>6ur>�2�>�}�>8�m    =��x>Ȯ�        =��>)I�>T�                 >�0                ?Cƿ?Es�>�                            L       parents[$l#L       #���                                                     	   	   
   
                                          L       right_children[$l#L       #               
         ����      ��������         ����������������   ����������������          "����������������������������L       split_conditions[$d#L       #@5��@�@@�n@
�1@"��'��@Q�?@4�=�Ո��&h@'��;F>�4���C?uY??묬��V�V�����=�04=Vg�ֺ�-���_=�L�?�J�� KZ?{/�=��:50k�Ԛ��:�=�G����;LAL       split_indices[$l#L       #                                                                                                                            L       
split_type[$U#L       #                                   L       sum_hessian[$d#L       #C��C�#�AwC��A"�W@~*}@�%�C�Z?���@�9�@�O+?Ƕ�@O@O]�@*�C핒?Ąa?���@=��?�>@�?�?��?�أ?�#[?ոC�<-A,�@^u�?�8C�F@�y�@8��@��@�-?��L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       35L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       O:�Q���|0=!�T<�q��sK>E�<�#d�+3>�[�l�h���[��>��*�u	�=��=w,�ax�>_�y� HW������ʉ�c�.=]�;8�=�\=���>��ʾ����>u�<�#��>L�/�Ո����V�e>��T���=�@Ǿ�Z�<ûV=���j�ξ�4	��
�>ǵܽ5��b�>�>����$pz��C�>����h>Fh��!�>�����>�|1�S�t>>�'�-�1>�����x����0���	>DC��԰s=BC�>�:�]�O?ջ<�J��<0<eR�<:˾�ڂ>̨�<��<L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       O                                        L       idI �L       left_children[$l#L       O               	                                    !   #   %   '   )   +   -   /   1����������������   3   5   7   9����   ;����   =��������   ?����   A����   C   E   G   I������������������������   K   M������������������������������������������������������������������������������������������������L       loss_changes[$d#L       O>A4r>���>)Yn>��>�B�>��>��c?*�>��>E�?��>-�=aq�=�>�>y��>�X�>�3�>�B>΀>��>!��>�Z?Sޱ>��>�T�                >6�~>Y9�>��?�    >�{�    >��X        =ɮ8    =�    >`*�>;�3>��<>��_                        >R��>PD                                                                                                L       parents[$l#L       O���                                                           	   	   
   
                                                                                                                 "   "   $   $   '   '   )   )   +   +   ,   ,   -   -   .   .   5   5   6   6L       right_children[$l#L       O               
                                     "   $   &   (   *   ,   .   0   2����������������   4   6   8   :����   <����   >��������   @����   B����   D   F   H   J������������������������   L   N������������������������������������������������������������������������������������������������L       split_conditions[$d#L       O�%Ʉ����A(�>:�f�%`��a�Z��D�Z�Ծ�v=�O��9v>��6�r
>��f��B�>�������̽�`g@��>�q?M#=�V�W���|��<��=� ���9R� gz�:`@�mw�2h�!�
�9,���׿G� ���	<��?��;��οC���>%8�ܹ,�V6>[�k��v5=:=ɏy�ESƻ��=�Y�@9�0@��B�=�
��<I=��o�~9Y=d�ɽPn;=�k�����m��?=k�ý�:$<i=2zF��.�># z;�X㽨H:;���;_<����=��?<C$L       split_indices[$l#L       O                                                                                                                                                                                                                                                                                            L       
split_type[$U#L       O                                                                               L       sum_hessian[$d#L       OCLT�B��:B�(B�%�BD�A5�NB�Z^B~�
AV�HA2�B0R@�`u@�\(@n�LB{ƈBV
�A"
A&t@CoP@��+@`�A�!A�@I��@!?��@��~@��?���@�ףBi��B/��A�5@�D@�a�?�.�Aǘ?̋X?�SH@���?���@��?��8@�¹@p�@�f�A�l@`>?��?��n?���?�|^@7�BT��@��B#!I@J�@)�@�S�@�D\@;+?���@���@���?��S?�9�?��K@���?��&@_�?��X@4=�?�N@�"dA���BO�e?�Ql?��@`0�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       79L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       59�=w����<�����uh�>��0<������g?���ē�>I*�;5��>>����< �����<v{�>�w�	<�3N�f�@>��X��dԽ=�#��.�U�D>��;��C>:�4��B��h�=mt`>ѓX�
?�>��,�S�=ݿ����)<�˾�~U�>C�>�$�=5
A��ƭ>�﮽'-���B�5�>�*8�#�>�j����L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       5                           L       idI �L       left_children[$l#L       5               	����      ����                  ����������������            !   #   %   '   )   +   -   /   1��������   3����������������������������������������������������������������������������L       loss_changes[$d#L       5>_L?ؕ?�q?l<�?@(]    >��?�    >�t�>UJ?Kw�?��?�~�?J                >�s�?0�j=� >ʆ�?�S>��?b�X>�9�?5�7?;j>��\>���        ?V�                                                                            L       parents[$l#L       5���                                               	   	   
   
                                                                                                   !   !L       right_children[$l#L       5               
����      ����                  ����������������             "   $   &   (   *   ,   .   0   2��������   4����������������������������������������������������������������������������L       split_conditions[$d#L       5>;�=��>T�D=��v?R��=��?�վ�#u>)�Y>Z>(�?z��?�C��;�=���.<;���=Ϣ���9?�	>�#z�k�N�H�J>�Ӭ@'�t=w�ʾ�k>>�-�?���)���<D=<�y=�}��]*�=�:��}D�<.!p�!�ƻ�n�;(�����dQ->I-<Y?���h=��H������:@n=�2��DA�=����MEL       split_indices[$l#L       5                                                                                                                                                                                               L       
split_type[$U#L       5                                                     L       sum_hessian[$d#L       5C�dCy�C;�Coc�A�\@J^�C8��Cm�?���@��<@�C*N�Af~�B0�)CAYE@�q�?�:?�_p?���CI"APWw@ީ@�TwB�|@�iC<�@�f�C�oAk:@�y@�u?��=@��@��?���AA�A�%v@��?�]GC:N�@#��?��@B�QB�31B�X@�2E@��.@l�@[��?�إ@�'L?��/@��wL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       53L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       �ax�9��վ�|3:�dI�f�V;I`!���9�������:��Q>��;��A��;:�l>A�&�g�y='eL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L                L       idI �L       left_children[$l#L             ����         	������������   ����      ����������������L       loss_changes[$d#L       >4N�>$>�    >6�;�� >n�s            >qT�    >,ۋ>B��                L       parents[$l#L       ���                                   	   	            L       right_children[$l#L             ����         
������������   ����      ����������������L       split_conditions[$d#L       @,�=?����>?�4���[�?�*F���޼�����?p]�=���?T�1�:`�=hx���(<Hk�L       split_indices[$l#L                                                                       L       
split_type[$U#L                        L       sum_hessian[$d#L       C��vC�&�?��C��@�C�M?�j�?��?�ZC�?���C�C$A(�C�NF@zoR@ް@fV�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       17L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       ?9Ќ)�/�`<���Xv༤�n<'
�>)S=S�n����>�V���i=;��Q�Z>�G��)>#}��n��hC���5��r=�� ��{X=�!��7��>HV��&3x��v����s>�Iq���d<�`q���>�Nd<�P��,>)�Ѿ���>|�߽s	�>�p'>⾳ߜ����=��H>g�W�oto>�c����w���+=�t,��=�X>�&x�éؾ;��>)o�S�<�?x�=�������<�|�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       ?                                L       idI �L       left_children[$l#L       ?               	            ����         ����   ����������������            !   #   %   '   )   +   -   /   1   3����   5   7   9   ;   =����������������������������������������������������������������������������������������������������L       loss_changes[$d#L       ?>@(~>���>d�)>�ю>�{>�Y3>є�=f�l<��    >�g�>�Z>���    >|m                >��?�1?� >��?B|K?&N=>#~->��R>�4~>�6>�>�?uP>� �    ?+bW?'Y�>m۔>�o�>m�<                                                                                                    L       parents[$l#L       ?���                                                           
   
                                                                                                   !   !   "   "   #   #   $   $   %   %L       right_children[$l#L       ?               
            ����         ����   ����������������             "   $   &   (   *   ,   .   0   2   4����   6   8   :   <   >����������������������������������������������������������������������������������������������������L       split_conditions[$d#L       ?��(�w��@�f����it�<�h�@,y���>do�>�W>ѯ����?o+s=�UT?�A=D/����Q������;�B�C!���͉�GϬ?�V@�>�J�?�N!?���=�|?��,�ԧҿ:Z�Kw<���(P�?R
?9�>?��,=�� ��Ү=ٹ�=6iܽ��"���<�FW=�-h���C=�μ�揽�H4=x� �i<�e�> }|���ѽa�=KR�~:;9؋> *t<�;��� �;�/L       split_indices[$l#L       ?                                                                                                                                                                                                                                    L       
split_type[$U#L       ?                                                               L       sum_hessian[$d#L       ?CI
�B��C �@�_�Bl��B��WA@!iR@��B?�:�Bh!�B���B8u)@P*^@��?�1�?��%@V]�?��B*u{Av�xBA�A�Y�B	�9A:��@9�@Y 
AՐB�@�&AlB<�?�R�A3��A���A��Ae?�Aw�@oo?��J?��}?���@��A��?�v.@~QqA� @�(?��P@w�@�>JA.�B%�A��@C�A=�AC�GAEu�@���?���AE��@�C?��L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       63L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       :��Ľ��.;�c�IC�>��>�>�;	�8����=�U>��C�#]��lI;�_���˘<��L>Yʙ:�\���{`�%��<�b>�?c��;���>���^w�>��;O�GL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L                     L       idI �L       left_children[$l#L                      	����      ����������������      ����      ����������������      ����������������L       loss_changes[$d#L       >9/\>�>��>G�T>�&�    >Y�	=�Đ                >D�'=��    =��>o��                ?6t�?�%                L       parents[$l#L       ���                                                                                L       right_children[$l#L                      
����      ����������������      ����      ����������������      ����������������L       split_conditions[$d#L       �Yt�<�UE�X �>Z&>�b�>�K�Rd�@�+<�f=㨷�D	;����E�?z�f<�a=N+ҿ#���-��F��<�;=�D�;n�!��=�޽�{)=��-:yJ�L       split_indices[$l#L                                                                                                        L       
split_type[$U#L                                  L       sum_hessian[$d#L       C�G
A,|�C��&A��@��?���C�)�@�M!?�rO?�ٌ?�d	@�C�!�@��?�jW@W� C�rx@�5?ǁ\?�W�?κfAfĉC�<T@�GAB�@��C�|L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       27L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       %��d7���9�;_����^=���|ݽ�Q���7=D�a���r�{51:đ�L��=7�-<�z2>�q�=�u⾝��>5׻��̻��b���>��]���=C�E���f>�Q�&���H_�䖅>���<U�b�p���>����	L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       %                   L       idI �L       left_children[$l#L       %      ����         	      ����   ����                  ����         !������������   #������������������������������������������������L       loss_changes[$d#L       %>��>��    > ]�>Q$�>���?0��>w��    >�~�    >�5�>��=���>/
I?MF�>.��    >p�h?�'?�~�            >PW�                                                L       parents[$l#L       %���                                               	   	                                                            L       right_children[$l#L       %      ����         
      ����   ����                  ����          "������������   $������������������������������������������������L       split_conditions[$d#L       %@,�=>]R��E��B�>���@r��/�A�̵v�
��V�` l��z�>��6�3S�)�>�]�<�v���>��0��)\������f=�u=��E�<j� �z�=�A��G�"�
��	'=�9޽{���w��=-ha�8�L       split_indices[$l#L       %                                                                                                                                   L       
split_type[$U#L       %                                     L       sum_hessian[$d#L       %C�ĽC��?��C��A��B��'C���A�)�?�|B��?��A+M�C�cK@���A5o6B�Y�@��?ʼ�A�:A\�(C�}r?ظ@W5�?�lHA%A�B�P@(�a@�S;?��@��@�RqA#ZI@e�|?��C��[@�Ŕ@���L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       37L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       /; �<^�D����<T�>��ž{�=}@�<O�P��%��_͈��ɽEY6>Z��:�}�=�u�=	�����>U���@��=�.\�r5�>��*��3�<@2�'�">���˕="�6��6�;�>������=w��x�>J~�;���>{�:>.�3�v���40O>6q�����>Ҹ�͸�<��+�������L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       /                        L       idI �L       left_children[$l#L       /            ����   	      ����                  ����            !������������   #   %   '   )����   +��������   -������������������������������������������������������������L       loss_changes[$d#L       />P>�>UԊ>@�M>)u    > J=���>-8    >RT>���>8ʥ=�z>���>i��    >#��=q�8=�y�=��            >i�.>��>k}�>J�    >3�        <�p                                                            L       parents[$l#L       /���                                               	   	   
   
                                                                                    L       right_children[$l#L       /            ����   
      ����                  ����             "������������   $   &   (   *����   ,��������   .������������������������������������������������������������L       split_conditions[$d#L       />��^>��?�wQ?��J=�S?���?�>?��ڽ��ƾ���?���>�ö?��?Ԑ�?c��<�տv�>Ο�>p��?�#
��Sa=ʝ ���?��Ⱦ���A�"=�<Cb�@�u;��=����V�z<������%=r��:�SU=�#=Qp>���]�X9�=Z�Z@=7cD����;�t��������!L       split_indices[$l#L       /                                                                                                                                                                          L       
split_type[$U#L       /                                               L       sum_hessian[$d#L       /CFzC/��A�|&C-�=?��A���@���C,߯?���AV'@��@q� @�C�A��?��u@�0@@!@��?@�&?�=�?���?�FWC�|AA� @MH]?���@��M?��?�"�@^1!?��?�<�?��tC}�@C.�?�R�@��W?�f�Aw�/@�o?�9�@�cw?��Z?�aC@��L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       47L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       a:�|ܼ��P<�%;����l�;�a�>jU='�뽏d�[{�= ���=_YE>�1\=oĸ�*L�=
1�L�G;�X��m���{~��f�>-�C<��J�W��>�?�<��>�'K=��y��&>��Ҿ��]�+�\��R�=�/���3���	���=��w���+>�����}>J��=nY���A>i�f�=B�="þ�$���?�=�P?�M���q��o>�*>6���E^�=�ݿ��R�j=���>1;���ї>���=��f����o{���>G�����<�ߌ>��<<��¿*z��o=���̈n>�X������F7)>�4⻲��>�&D�:o���5�eN>�w=�Y??�O���>K^�>��z����W�9>�������> ;,L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       a                                                 L       idI �L       left_children[$l#L       a               	                                    !   #   %   '   )   +   -   /   1   3   5��������   7����   9   ;   =   ?   A   C   E   G   I����   K   M��������   O����   Q����   S   U   W����   Y   [   ]   _����������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       a>7%d?	ss>��S>���?4\>��t>��v?�v? Y�?�KC?[�?��?� .=$�>졞>=J�?m\?LdW?W԰?[�>�>��}>�!?K0�?=n>��>���        >퇒    >{��>%Vd? 6?v�>>`�X?o>��>���>��    ?:ϖ?C�        >zz�    ?��X    ?��?��?2�*    ?�?�L>��9>��                                                                                                                                                                L       parents[$l#L       a���                                                           	   	   
   
                                                                                                                       !   !   "   "   #   #   $   $   %   %   &   &   '   '   )   )   *   *   -   -   /   /   1   1   2   2   3   3   5   5   6   6   7   7   8   8L       right_children[$l#L       a               
                                     "   $   &   (   *   ,   .   0   2   4   6��������   8����   :   <   >   @   B   D   F   H   J����   L   N��������   P����   R����   T   V   X����   Z   \   ^   `����������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       a������5�?�վ?h͆>�2˿��?βH����?���>�Ӭ��e �?�a��t��V�2��>�"U�e��?�zn?���
��,��?u(X�� ?+1�>�Ӭ?QZ>}�=#I�]*�=�斿hy�>�ŵ��z���k�����@�D�д?��?O��=�.���?��J<���	����Fʽc��M@�I-?��2?�~[>�����U?�U��"��F�@
k�<�����彌g�=	��=T�۽�>��<�cH��t��Ǿ
u�=5����6<�>�$<	�u�1̓����=�@��p�=��⽲9)�m��=�?v��T6=�ǅ�_�+�*@�;��>Gy<�h�>f_��(=t:=��,�yA���#=إ����=@GL       split_indices[$l#L       a                                                                                                                                                                                                                                                                                                                                                            L       
split_type[$U#L       a                                                                                                 L       sum_hessian[$d#L       aC�7(CM�Cb�IC!a�B2#CO-�A��B� BD0�A� A�&B��"B�hp@��AfQ*A@BB��A�A�A� ]AD��Ak�@��$AO/:B�v<A��@���B���@g$t?���A<>Y@(KD@�M@�|6A���B�I�@��A.�@�(A�_A4͊?��A{D@�.�?�7�@?8TA6ۏ?VB�m@#�A��@�@��?�8HBw�Aߣ$@�o@��?�k@��?��@H��Ab�Aek@�ElB�e�?�@��@(��A�B@@ �?��c@F�A�6>A�@+A@��@��@h��?�E�@T�+A��B���A-��A|߹@���@<��@~I@!��@X9�BYo�@��AR��Al�n?��@^�-@���?�_kL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       97L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       -� ��;"潗8���eH>p夻��ᾊ�9_z�����>�����0F=L�#��`���q��E�;�+��n���@?���b&>1'N���d>b��qyd��a¾X>*>N�~;r>�v���g��7r�|>#�|c>g<;����=�T���=�2�#A�=.�(�q7>����`�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       -                       L       idI �L       left_children[$l#L       -               	         ����               ����      ����������������      !����������������   #����   %   '   )��������   +����������������������������������������L       loss_changes[$d#L       ->|S>�a>�Ef>y�Z>���>�po>��4>C�    >��>8m>�$�<��`>L    >���>�                >�>�/�                >�6    >i.4>��F>�        >|x                                        L       parents[$l#L       -���                                                     	   	   
   
                                                                     "   "L       right_children[$l#L       -               
         ����               ����      ����������������       "����������������   $����   &   (   *��������   ,����������������������������������������L       split_conditions[$d#L       -?-M�?������?^h>�9C��tB�Ž�?�G���*0��?&��=�6���dy?�.B���S?��Ⱦ"Nv�ـ>�����=T���Q�>2$���p��uP����=w��?��Q=����>	D?HO�=D�ѽ�4	� ^�:��a�
7<�q ����=��C�6<Q�d���!=�"d���;L       split_indices[$l#L       -                                                                                                                                                                       L       
split_type[$U#L       -                                             L       sum_hessian[$d#L       -C�#C�vzAٺ�C�)�@�+�A�I|@��nC���?�C#@|g@)�.A�d�@7'1@,�
@^��C��Ar{�?�0@1�k?�Z�?���@��zA%Io?��?�]?��?���C�M�?��M@��A+@�*+?�U9?�JA -C���?��p?��6@[j�@�G�@��S@o�@��P@�2�?�7JL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       45L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       S:�]꼵�=#��<s�h���6> {`<��p�(�>p�e�Խ�<g�>�^C�P=/�<�(��[4;M��>�w����Ѽ��7�ZM�<��g���>�x��Ln=�m>��
<��p>����C��{[���>X�8�k�>�{ʽ�)���<�r�=��kO���	9���>�"+��Z�hɢ=�JF>r.��W�=��q>�('�J�=�����'?B����8=9��H��> YѼ؁p>��<>�X���\���t������>?8����~;Ec>F�g��
>�f9;Ip�r5|<���ZB���S=�R�>�X�<����\��<�2�>j�vL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       S                                          L       idI �L       left_children[$l#L       S               	                     ����               !   #   %   '   )   +   -   /��������   1   3   5   7����   9   ;   =��������   ?����   A����   C   E   G   I   K����   M������������   O   Q������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       S>8�>���>>>_9>�΁>���>]�?[q>� �>#
�>�2�>Va�    >p�>[L >J|>��*>�"5>� >�h>
W>5�?��>
�:>%�        ;�@>EC'?i��?X�    >�{>l�>ݎA        =y�p    = H�    >4>�>]}�>m<�=FV�    =K�            >���>a��                                                                                                                        L       parents[$l#L       S���                                                           	   	   
   
                                                                                                                 !   !   "   "   %   %   '   '   )   )   *   *   +   +   ,   ,   -   -   /   /   3   3   4   4L       right_children[$l#L       S               
                     ����                "   $   &   (   *   ,   .   0��������   2   4   6   8����   :   <   >��������   @����   B����   D   F   H   J   L����   N������������   P   R������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       S�%Ʉ������>:�f�%`��?���m��Z��>C��=�O��9v>��6=�
�?O��B�{;�">�Q��C@��>�q?M#=�V�=^��;f���(�=�>6$�?		��E�D�f�K�}7�9,���>p��>��-�2?��;�VH�C��/�=;F]��bC�V6>[�k>�8�<��m����<�"=Ȗ��P ?2R�4�/>�l��̪<^�ܽp��=@kȼ�D=�q|=����7�� ��B��
��=ew'���1:l�;=nK��28>��:#�T��SK;7����9��e�<�0=�jv;��ʽ�cS;��F=�خL       split_indices[$l#L       S                                                                                                                                                                                                                                                                                                            L       
split_type[$U#L       S                                                                                   L       sum_hessian[$d#L       SCC��B�8B��B���B:-AldBn�>Bw�PAMPA"�SBnEA#��@�.C@K-�Bb_BQ�AH�@�k�@�4|@�A(@Uj�A��A��@��7@��@t|?�r�@)�BWj�A=�B"J�@F�@�nv@6X�@�?F@K�x?� @���?�`�@#B?��r@�	�@i+�@���A��@B�M@ �"@V�K?�%?��?��!A�kyA�i�AX�@Z?@��.B��@��8@�|?��W?��D?�=q@w��@�I?�X?�s�?���@��?��?��3@'�e@2�V?�_ @po�A���@ ٠?�OY?�1{?�EAȰ=@���Ax��@��L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       83L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       5:��V�-F=�,��=k����<���>U@������O�=Ө��>Ҿ�;Ƒ��FB<�{]>��=P2G>v�὜�>����� �R�><Z��� ż��e>�Iþ�(=�L<�(>���=`j��r����> Tż������G=�H�?H"����<����3��{����>+>L�ž������$>��=���N���=ɽ�@�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       5                           L       idI �L       left_children[$l#L       5            ����   	   ����         ����                     ����   !   #����   %   '��������   )   +   -����   /   1   3����������������������������������������������������������������������������L       loss_changes[$d#L       5>.�>�b�>���>�"�    >�<>��?    >�,
?�N?4�    >��?F��?2^�>��L?��>���>ƴ�    >���>炁    ?`�?��`        =���>�>���    ?Z��?.7�<�                                                                            L       parents[$l#L       5���                                               	   	   
   
                                                                                                     !   !L       right_children[$l#L       5            ����   
   ����         ����                      ����   "   $����   &   (��������   *   ,   .����   0   2   4����������������������������������������������������������������������������L       split_conditions[$d#L       5?0\�?.�?��b�Ծ��<�5�?�C����;�P�YQ���:m=��?�S��N���DZ�]��U�'�?���=�?�(X��B��(c���:��$��˭>,B�V�|�(��?�i�>	��?k8�?tt�.�"=@e����潶c"=�->7�)��B=;��o�����J����=M:q=uú�� ����>�	<艠�wBf��J%�&�L       split_indices[$l#L       5                                                                                                                                                                                                 L       
split_type[$U#L       5                                                     L       sum_hessian[$d#L       5C��C���B���C���?ھ�B̾�A	��@9YC�PFB ��Bx�0@q��@��TB��CP��@���B-@�i�B\��?�@`��B�J@o�A�ǣC:��?��@~2�@�MB�8@}�'@B�Ay��BQ@�?��9B�غ@�Y	A���?�@ꉢC3ff?���?���A$mA��:@3Ҥ?�AA/@c6�A��A��=?�q?�[�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       53L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       ;��̸:kWV��<��[�t>=�5h=��U��6�>ݩ�퇥� Ɋ���<��|+;���A��>��)=8����<> �S7�=f�=��6RU��-�<��?.��
C><��
3���徝#,?�<�$ۺx���l�>W틾 �_;��P>>�н��t>H��]��݈>Xc6�7{Q>k�s?-�,�uZ�<��{>��M��;ܢ~=���h��:�93=�<��/�>!,����L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       ;                              L       idI �L       left_children[$l#L       ;               	   ����      ����      ����                     !   #   %   '   )   +   -   /   1   3   5   7����   9��������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       ;>��>��>(y? ]?_�=�'     >���?]N�    >�*�>�-    >��>��??��T?E�H?JU�?��=���>'��?a�?^;� >sb�=dn�=V�?,�?�i>��
>�\h    ?                                                                                                        L       parents[$l#L       ;���                                                     
   
                                                                                                                          L       right_children[$l#L       ;               
   ����      ����      ����                      "   $   &   (   *   ,   .   0   2   4   6   8����   :��������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       ;?
ڿ.p>����&0��_¾V�<�O��-�d� �o���?�ͨ<�0���g>�� ?��b?{/�>fނ?EU	?�	L�9��rI>��?V��DFZ@c�%J�?�>�Y?`��(������>70�3���No����=����A0:�Xa=d���ь%=/;����=
=��!�\-�=�x�>P���6�;���=����8���a=�"���09�=���/=AP5�ň�L       split_indices[$l#L       ;                                                                                                                                                                                                                        L       
split_type[$U#L       ;                                                           L       sum_hessian[$d#L       ;C��C�0A � C_5>Cu�!AN?�N�C:8�B�?ߩ\Ct�@���@ .C1܅A��@���A�bCg��AB�!@7�/@=:�Bޅ�B�3u@��	@��@�2H@�yA��AI�C_�HAHG?�=A-�:?���?��?�H-?�-�B���A�OB\��A7l�?�7P@A�j@��@�+?�M@�I�?�~Z?�AG#�@{�;@��b@��@ʜ�CY�c?�ES@ο:AG`@!�gL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       59L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       ;�t;��־;-k>U�q;'/J��x�=.��=2nG>�r[����<!/���艾�9<>��;G: ��6<N��>2����L>���;�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L                  L       idI �L       left_children[$l#L                      	����������������      ������������         ����������������L       loss_changes[$d#L       >'�o>�)>50�=G[�>��                =S��>�d            >t�T>�8>��j                L       parents[$l#L       ���                                   	   	   
   
                  L       right_children[$l#L                      
����������������      ������������         ����������������L       split_conditions[$d#L       ?:h��p�e?�C=�+��o�|���M<Q�<V�=�V��겿nY�����w�=ȃͿaD@�|���`Q�=����E�=�F;e�L       split_indices[$l#L                                                                                      L       
split_type[$U#L                            L       sum_hessian[$d#L       C@��C<�@k��@+ 8C:=�?�D�?�Ϊ?Ȱ?�Pc@V�C6�?��=?��@6�BC4TA/]#C)�@bO�@�M?�	#C'�oL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       21L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       %:��q�W��=�@~:��¾��6>�)<�}?��>�b�=�N��%���>K��9�&���9�>h��������}>���By�;��H����>پ���d=N�o�e��>VK�8�9���ţ>�2h:�bӾas�>�;+����<� �=�Id>�EL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       %                   L       idI �L       left_children[$l#L       %               	����      ������������         ����         ����      ������������      !   #����������������������������������������L       loss_changes[$d#L       %>Gi�?��?h5?��?Iv    ?p'>��            ?(^?#>��P    >�:N>��,>��n    >�,y?9M            >�+�=ы�:�-                                         L       parents[$l#L       %���                                                                                                              L       right_children[$l#L       %               
����      ������������         ����         ����      ������������       "   $����������������������������������������L       split_conditions[$d#L       %?�p�?���?�?�?ڈ?A�[>��zz?�mO>$=bs�,�6�O<�>v�,�g�i�	�?5@�澀lM>	P߿r�l�e���X_>����p�>ec=�k��'7�xʾ��>Qr9�˽�E�=�ν�Y;��<�$�=��zL       split_indices[$l#L       %                                                                                                                                   L       
split_type[$U#L       %                                     L       sum_hessian[$d#L       %C�_C� @A��(C��*@�P@2!aA���C��X?��'?�WH@&^�A��A�C�+5?�"�@)�@�^@�4�@\�	A��C���?��?��}@�1�@��@'�Z@��@�'�@Ik�?���C��?�)�?�p(?�v?��>?���?���L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       37L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       5�y�;P���5f�#�>�Ft�~���	:v,~��;ٽ#�>��c="Ͽ���>ɨ��g%�HR>by^��9'���H�4��=�rq?5˜>^%�M�[>޶�=#A?�N=��R�?�V<Â���Fx>���u|�=�82��P�����>�b>�׾��M����>�p���L��D~��ɾ>{�y�����=>=;I�Q�U>�
=��o>YQU���OL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       5                           L       idI �L       left_children[$l#L       5               	                     ����               !����������������   #   %������������   '   )   +   -��������������������������������   /   1����   3����������������������������������������L       loss_changes[$d#L       5>"��?@LA>ƫ>�2C>���?/ ?��>���=�@=��f>4E�?��    >^DL?Z�>M�;?^�>2�	                >�Y>>���            ?W�;>�Q4?}7�?n��                                >�A�=�Y(    ?F �                                        L       parents[$l#L       5���                                                           	   	   
   
                                                                           '   '   (   (   *   *L       right_children[$l#L       5               
                     ����                "����������������   $   &������������   (   *   ,   .��������������������������������   0   2����   4����������������������������������������L       split_conditions[$d#L       5?΄?� ?묬?���?e�m�)
3?�ۑ?�Ę>�ŵ?�4P?�۸�"(������7?��D�k=	���s|��W�Y_=w�>Z'�?�k~?
C>��<5]�>5&^?5�J�-��[��ٶ>Z��J�=
!����#��>�=(�6�Q�@�?��J�͔�#v���?=����˒��=c�{�g>lg<��=�d ��#,L       split_indices[$l#L       5                                                                                                                                                                                              L       
split_type[$U#L       5                                                     L       sum_hessian[$d#L       5C�'C�vB��C���@�U�@��A���Cӑ�@���@"^�@�&@_��@��@��A��C�#�@�{�@1*�@]	?���?�?�!�@A;B@��?� �?�u�?��AeYSA]�mC-2ICu%@>��?�
?�x{?��&?�[?�j?��_?���Ao&@��Y@L-A*��C3xA���A9�Cl!�@)��@��@A>E?���@��k@��XL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       53L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       G:�S'����=6E<Auw����<�>8yC��f^=��2�/�l�`�p=(��,�C>�-�<ǥ,;�C��cl�>�ޫ=M�S�i���?�⾐5J=}�<��>��=Vt۾�ɕ>I�$�xC���W>�e�F���ʱ�L�M=�>���J%=�>�4���#��9;N%�=��M2��V&�>�Ӗ>~u�,�"='4�>�k<rM+�%Ž�n>���>7�Ǿ��8��C<�м=�>s�b���=��y��qh�)<}n>�|#=�a����=��p����>���OpL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       G                                    L       idI �L       left_children[$l#L       G               	                        ����         ����   !   #   %   '����   )   +   -����   /����   1   3����   5   7   9������������   ;   =����   ?   A   C   E��������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       G>�>tQ>	)(>G��>]�~>B	>5�>���>\>H{8>2�v>"�<>u"�    >�<�>�'�=�h    >x�"=�`h>>{�>5d    >�cV?ٰ>8�	    <��0    >9��>{�    >���=�w(>�            ><9�=��P    >�f4>:մ>mr�?2�                                                                                                        L       parents[$l#L       G���                                                           	   	   
   
                                                                                                     !   !   "   "   &   &   '   '   )   )   *   *   +   +   ,   ,L       right_children[$l#L       G               
                        ����          ����   "   $   &   (����   *   ,   .����   0����   2   4����   6   8   :������������   <   >����   @   B   D   F��������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       G�K�l�-��@�|�j�;*�?�U�@�ھ���i+Y�4?�B?��?���=��?�j�?[/D��=�q��J��?1d�ݑ�?��`<��?P��?X<h�����XM?�>Խ����Q�H�0���!������� g=Х*�¿`<#̯=�r~@	�F@ª:w`�?gѾo��?��v?c��=����O<)<H�~=���;�a��&� �:�Q=�4�=\;V���D���
;�`�<=��=�Vn����<��žD�)Qe;��=�a�<�tv��|\<�����"><��xt!L       split_indices[$l#L       G                                                                                                                                                                                                                                                                       L       
split_type[$U#L       G                                                                       L       sum_hessian[$d#L       GC?��B��B��SB��B%[�B��@��B\�KA���BTeA �B�"�@r�?�ʶ@\��BG@�b?�A�ݔ@y;�A�S@��F?��B]��A'�@W�?�];@7n?��B9�0@S��@c@Ha@B�A��8@/�U?���?���A��@�DE?ִBL��@���@V�@�#�?�F�?�i?�Z�?�*Bn$A�.?��y@\�?��t?��?���?� *A[�}@w��A���@߸W@s�?��B@��@A�h?���@<�C?���?���@}�@,�CL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       71L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       #:����V��=��:���R>��<��y�'��>ݺ,=�]:�����1�>L���ռ7�в�ҖǾ��˽���>��A�/�8;��M��0>7_پ���>1��=��V>�|��S6<���?�9:|���[��ޘƼ��>�DL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       #                  L       idI �L       left_children[$l#L       #               	����      ������������         ����   ����                  !������������������������������������������������L       loss_changes[$d#L       #>2�l>��>��?	�>�^�    >隟>��            >ⅴ?��>�u{    ?+�{    >�1=
��>ҏ�?E�|=f�@>�	B                                                L       parents[$l#L       #���                                                                                                        L       right_children[$l#L       #               
����      ������������         ����   ����                   "������������������������������������������������L       split_conditions[$d#L       #?�p�?���?�?�?ڈ?A�[>��?*~V?�mO>	N<��F�p�?$��>]G�g���oQ�1����@
6?) �>��P�e��B�f=D�����=U�=K>A���u;���><O�9�7ϼ����޻��Y=�Q�L       split_indices[$l#L       #                                                                                                                            L       
split_type[$U#L       #                                   L       sum_hessian[$d#L       #C���C�<A�gC���@��@!t0A�8�C��7?�?؇h@%��A!��@嶬C�N�?��A��?�_�@S��@w�qA�cC��@2��@�ņ?�C�?�TE?���@6�@i��@�w�?��pC�_�?��j?�; @]��@ˌL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       35L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       '���:�����o����>��s=F\u��]�:ͭ'��C�<2��?:a��8>CA�=6@���Rǻ#b�>z��P��>aቼqW?���&>����!.�?Q�>�%:�+�~������>��G>��g�o7>�]!���!�;�>�3����=��>ޜW=L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       '                    L       idI �L       left_children[$l#L       '               	         ����   ����         ����      ����������������      ��������   !   #����   %����������������������������������������L       loss_changes[$d#L       '>�^>��g>�f?!�>��u?�}>��r>�n    >J�    >�>���>�o�    >��?�                >���?6��        ?�>��l    =�w�                                        L       parents[$l#L       '���                                                     	   	                                                            L       right_children[$l#L       '               
         ����   ����         ����      ����������������       ��������   "   $����   &����������������������������������������L       split_conditions[$d#L       '?�p�?��ؿzz?ڈ=3��O<��U��?ͩh��'?�b�>-�?5?��(�V�z�1�?Ş�Zo��z[�=��S�����H�?+�;�L���e�A=��?�(%������P>�ؼ��j=�<������?p>���q[=��>�<>��L       split_indices[$l#L       '                                                                                                                                            L       
split_type[$U#L       '                                       L       sum_hessian[$d#L       'C�gC��A�8C�.d@pA.A)L�@�GC�D�?�o�@��?�T@D$@�~@;[@���C�`@˥?��B?���?���?��@�G�@8��?���?�.AC���@�L?��@�+@H�f?�r+?�??���C��?�A{@VE?���@��p?�ʣL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       39L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       :hB;Ǖ�/�;ߣ>�/��WK> =<&h��ßZ��o���V;��7>��!�,^�=ۋ𽤫-���D<&2�E�\=q�9�^�D��F�>m��;�}�>�I������뾏��=��<L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L                      L       idI �L       left_children[$l#L                   ����   	����         ����   ����      ��������      ����   ��������������������������������L       loss_changes[$d#L       >�`>4 ,>�>J`    =<p    >1��>c�d=>}    >�M    >W> h        >���<��    >4L                                L       parents[$l#L       ���                                               	   	                                    L       right_children[$l#L                   ����   
����         ����   ����      ��������      ����   ��������������������������������L       split_conditions[$d#L       ?���?��@�R>��^=�>p��=2J>��?�B��q!��>G�=�������?Q���Ś7�ё�=��Z>���<�$�@�u�ڻ�=��:�c�=�X|��L��=3���N;<�B�L       split_indices[$l#L                                                                                                               L       
split_type[$U#L                                    L       sum_hessian[$d#L       C=�C7��@�+C5��?�dX@��?�E�C(�#AM\�@s��?�-8C'n]?�c.A7@Q�?�r�?��\C%'�@�K?�z�@�ϸ?��z?�^�C"��@�K?�w�?�ȣ@�ܽ?���L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       29L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       :��)��0 ;����J�>w�>őh;,�꾬�ֽCqd>���Є�~�[;��Z�
a>��>lWs;2D��j``=���ĺ=:k��� ;Ѥ�>�e�<��L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L                    L       idI �L       left_children[$l#L                      	����   ����   ������������      ��������   ��������      ����������������L       loss_changes[$d#L       >3uL>n�L>�W>.�$>r    >>r    =��            >!R=ʿ�        >%��        ?��>�M�                L       parents[$l#L       ���                                                                          L       right_children[$l#L                      
����   ����   ������������      ��������   ��������      ����������������L       split_conditions[$d#L       �Yt�<�UE�X �>��P>�b�=��Rd���ih����=��i�9���ޝ�J�T>���=9�2=��?0�r���:<� �<�h�?F#\��4:���=��;�NL       split_indices[$l#L                                                                                                  L       
split_type[$U#L                                L       sum_hessian[$d#L       C�4?A�)C�6m@��F@&?��Cʆ�@[��@��?�f?��?��Cɐ�@Q�?�'@��CȊ�@�?���C�
�B� XBhWC�}�@�ϐB�c_L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       25L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       E��ޏ=#r4����P��>��̾�xh��7
=�J�\���d>��s=�O���-;e�N��3�>11q����>z?�)>+�`�%�˾R�e����>>	C��E	e��kT��� >��U�JƑ>#Q��Ҿ!�g>���?�?>�X>���Eþ�~;����>����	��%�>������L:�t�*1�>��{>��b=�!O��̱>�v����>�BQ�����0�>C�羗G�>LG�HR��F=���>͌	�:���K���->����/�'L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       E                                   L       idI �L       left_children[$l#L       E               	            ����   ����                     !   #   %��������   '   )   +   -   /����   1   3   5   7��������������������   9����   ;��������   =   ?   A   C����������������������������������������������������������������������������������������L       loss_changes[$d#L       E>	�?�λ?�=�?$.?b�J?:<�>��>>�2_?Md    >_:�    <�# >���>���>���?�?��g>�
�=]=�>�4~        >���=�1 >��>�0>� M    >sX�?)��>)�>8��                    >p�x    >9J�        ?�_>���="�P>QU�                                                                                        L       parents[$l#L       E���                                                           
   
                                                                                                                 &   &   (   (   +   +   ,   ,   -   -   .   .L       right_children[$l#L       E               
            ����   ����                      "   $   &��������   (   *   ,   .   0����   2   4   6   8��������������������   :����   <��������   >   @   B   D����������������������������������������������������������������������������������������L       split_conditions[$d#L       E�[���]mZ�Z��`ن�(h�\������f�* 콚��09�=
�q>���>/@1�`���f�f?2��>AA�`)�?jN>��P�F�'�|�����C��)r�Vix�gt���.g�c'�>��(�_AK� PͽBb=��>:��=+rj=��}�J5���dG?__=���9�+�>�Ӭ��`g�T���L;n=��=�<��ƾk=�n(��Ǎ=�O��)�SYU=j�����H=u#�pb��Ü<�J=���_;=�����j=��ȹR�/L       split_indices[$l#L       E                                                                                                                                                                                                                                                           L       
split_type[$U#L       E                                                                     L       sum_hessian[$d#L       EC�S�B���C�,�Bwy?A' �@��C��%BI,uA93'?�N�A��?Ѭ{@���A#��C��FB	a�A*�@�ސ@qz@�#@U/1@oJ�?�h@�W�@E�(A���C�'�Bv�?�[uAP�@8��@&@�ˆ?�,@��@��?��?�a%@��@��N@+d�?�#%?�]*A�HA*@��C��A�"�@&[W@�_Q@���?�Q�?�r?��?�g�?�a@��?���?�Vv?���?�4?���@��@��Q@!��@�@GN?�^�C��L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       69L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       A9�$���8<��<�O���t���=���G�r>�{���4�KU< ��n�o>x�B<���>���|�>��Z��\���jؼ�)�����>ljt�������>���w��=,�!�d�>��;�^P���:>@Z���J�=�HH�2<���<d�Ӿ�4�=�v�>�I1�*�6>1��<���>��z�OR*>5�¾�wܼ�u=���Bq�>��I�o{�s��=Q	�����<A�=��L�>,�$>�%H=�莾�=�s<>�FȾY]L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       A                                 L       idI �L       left_children[$l#L       A               	            ����                     ����   !����   #   %������������   '����   )����   +   -   /������������   1   3   5   7   9   ;   =   ?����������������������������������������������������������������������������������������L       loss_changes[$d#L       A>\M>+��>Þ>�W�>~0>�^9>��*?My�>�G    >Oy >L�B=��L>2�l>GC�>]Y�>���    =�P    >k�g>�z\            =��x    >xM>    >Z`>�Q=�&x            >#ۘ? �b>@_2>$��=�=���>�_??�R                                                                                        L       parents[$l#L       A���                                                           
   
                                                                                       #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *L       right_children[$l#L       A               
            ����                      ����   "����   $   &������������   (����   *����   ,   .   0������������   2   4   6   8   :   <   >   @����������������������������������������������������������������������������������������L       split_conditions[$d#L       A��8�/)-�1��>�x�2V��à�QB������I�Ő��*p.@䲾?���@BN���?-B=�e����Ҁ7=���?� j=��y��Z�"��%[����V?		���X��h\�HM^��nD=f�I���<��$�1�><��29D?�i�z>̎�?M�?�;�i�>X�x� =ZV��؏ջ��<�:�iUW=��X�6�.��,�<z�Y��D/;ho}��\==O�>��<��޽B}<�W=��k	L       split_indices[$l#L       A                                                                                                                                                                                                                                            L       
split_type[$U#L       A                                                                 L       sum_hessian[$d#L       AC<"�B��0B�UA̢"B$�PB���B0#�A�@�pZ@0;%B�B�!@n�AqBb
A&[ZA��@Xw@�=?�Q�B�B�}�@3��@%��?��@�xT?�R6BbS?���@��@���A�?���?���?��A5��A�):B�ƃ@v��@`~@�HAƌ/Ap�@ �k@D,@(��@X�@�j�?�2	?��|A��@(��A�!A���B2��@��?��?�2�?��B@V��?�҈A!9<Ak�"@�*�?���L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       65L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       :�G�
�;{4==���̶�>k'�9��!��>±�>�𰽉�Y��(�:Ɗɾq[}=����0A?2�־���>��>�~}��%^��/E���a�j�f;Q97��md>4��>��-8���L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L                      L       idI �L       left_children[$l#L                   ����   	      ����      ����   ����������������   ��������   ��������      ����������������L       loss_changes[$d#L       >,*>�F�>�ފ>��?    ?9n>�.z=���    ?��>�Y�    >�>�                =�|        >�        ?xd>�Z�                L       parents[$l#L       ���                                               	   	   
   
                              L       right_children[$l#L                   ����   
      ����      ����   ����������������   ��������   ��������      ����������������L       split_conditions[$d#L       �j���l���g�D�m����>��f�f?:=��7�6?P�l���t�fｐ�<����9�>V�ν�^=�BS>�c����S��u�PI��b����=X� =���7�&�L       split_indices[$l#L                                                                                                                     L       
split_type[$U#L                                    L       sum_hessian[$d#L       Cή4@ߩ�C�/�@�%@/l@���Cǫ�@G�
?���@r(�@O�f?�qYCư9@�e?�}K?�n�@qw@5,?�&t?�f�C�	�?�,!?�>7@�pvC��@�R�?�v @$�C���L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       29L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       9����:��
���\;�x�nT�>�>�)�:��6>���u�b��3p>_uJ�q�ξ|>	�i��;�[�o>>�Ӯ���%<�%����~>��ýU�o��#ɾ��}>�]��S;�>UK��eI���P?� >T�8�6?�>��u=�O?�(=��e�,yӾ�q𽍧c���<<ٱ��>Ԫ>�WZ�e�+=��c���6�'�>��=�9E������[>��X�ڃ⽃X/L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       9                             L       idI �L       left_children[$l#L       9               	                  ��������               ����   !����   #   %����   '����   )   +   -   /��������   1   3������������   5   7������������������������������������������������������������������������L       loss_changes[$d#L       9>��>�F>]�?$�7>�x=��=���>��\>Ҷz>�&�? d        =UP=��g>r�=��D=é�    >�-g    ><hz>�J!    = �    =��>j�?>1n>�4        >�?�>Z��            ?-n!>���                                                                        L       parents[$l#L       9���                                                           	   	   
   
                                                                                         !   !   %   %   &   &L       right_children[$l#L       9               
                  ��������                ����   "����   $   &����   (����   *   ,   .   0��������   2   4������������   6   8������������������������������������������������������������������������L       split_conditions[$d#L       9?� ?΄�h�?� ?묬?���?�7�?���=�C�)
3?�ۑ=�-���⾆��@ټ?�Ę>�ŵ?����kǿ0���/L��7?��D��^%?�5=-�p=��a?���=	���s|��=->7	�?ʿ&�2�=�&<+#,>'h�?5�J�-���U�������<��4�L="�3>4j��д=�o��	۽� >
P�=�������;=�NѾ�L       split_indices[$l#L       9                                                                                                                                                                                                              L       
split_type[$U#L       9                                                         L       sum_hessian[$d#L       9C��7C��	A?��CϠqB��@	��Az�C�?�@��@�EA遫?�~N?���@�b@��JC��@���@��W?�Va@T��@x��@c�A�52?��y@B��?�R@h�kCǮ�@��@+��?�eM?�C@I� @٣?��V?�+|?��AZ�$AQ�@?��?��k?� ?��C�w@���@5�!?�	?��R?��?��Z?�Q�?�pr?�B�A�v@��]@8t�A#�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       57L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       G9�(<�IZ��l�<��9>@�-����=� <�6�F��>������^�$s����=�2��U�;�G/=��<��龎�>�-�=�I
�:�A=�G>�>߽Fj>�[���n�8��>Ѿ<��5�U>�Ju<F���S��=}=���8���3�>�o;�;ɾ��>Ua���y>�>�>��;е�>u�S���i;�l�=�<�>�D��k�M=�����P�0>tf�I�>ٞs<��x��9�>�+ܾ���=}>�j���>!�߾���>���=<I�>a���_L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       G                                    L       idI �L       left_children[$l#L       G               	               ����                  ����������������   !��������   #   %   '   )   +   -   /   1   3   5��������   7   9   ;   =   ?   A����   C   E��������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       G>�c>(~�>�v>=Q�>f�>yZ�>#+H>т=�.= �    =��>�7�>� 3>��C>X�>�/w                =�3P        >|J >F�>��>�@5>�p�>_�V=��@>+)�>W�=        >7)i>.x>��>�4�>�O>�Bj    >y�>�B�                                                                                                        L       parents[$l#L       G���                                                           	   	                                                                                                     !   !   $   $   %   %   &   &   '   '   (   (   )   )   +   +   ,   ,L       right_children[$l#L       G               
               ����                   ����������������   "��������   $   &   (   *   ,   .   0   2   4   6��������   8   :   <   >   @   B����   D   F��������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       G�d�?K�?\Kb>�\���~=��E?���|�j�/
 >�����@'�>𰽩��?8L��=ץ�;�>���c�=�j<��@�k<�S�=�?��e?��@A>�~�:?�T�?[/D�� g�>:�f���D<��ٽ����v��N��?�i�>���>!W��G�8=:�7�V?���:�s�=������:���=	��>)?��O�<��L����1�M=4���r%�>�E;�����=��<��A<���=���1�=B=s����>k�<a�?=�_Z�흦L       split_indices[$l#L       G                                                                                                                                                                                                                                                                  L       
split_type[$U#L       G                                                                       L       sum_hessian[$d#L       GC9�rB���B���B�U�@���Bp��B^7B�u�@;��@p��?��A���B)PLA��MA��!B���A}�^?��?�D�@,:�?��A���?�f�?��4B#Y
A��AH�A��@���BphP@�Ȭ@��7A-�BAs�?���@3*8B&f@�t�@5)@�b�@���@��?�k�@�@/ߣBc,@S�@;��?�a@]��?��!?�;A�;@,��AG�<@�S�B��@�}L?��?���?��[@m��@c6�?���@ň?�;1@��@�i@m�?�Ź?���L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       71L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       /:��ͻR�=��L�1��:i2>i3<�
����!�#?�(�Ͻ#$Q>���>0ѽ��%��X��ݙ>��ؾt�K;�k�!L=Z�>��k�|`]>�&��v�=醼����=��"9�t>�.�>$�g��4�>@/��EV��S��
�a>���t���^�<R��n>��H����>'V">��8�*�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       /                        L       idI �L       left_children[$l#L       /               	            ����   ����         ������������         ��������   !����   #   %��������   '����   )   +��������������������   -��������������������������������L       loss_changes[$d#L       />�?>�k�>*�A>o�? �S>*p>X!d>��?�    >��X    =t��>���>�v�            >VK�>���>�#8        >wHL    >GH> r        >wAf    =�{[>�B�                    >�;                                L       parents[$l#L       /���                                                           
   
                                                                             &   &L       right_children[$l#L       /               
            ����   ����         ������������          ��������   "����   $   &��������   (����   *   ,��������������������   .��������������������������������L       split_conditions[$d#L       /?ܭ��g�@SM>��P�e�@�\_�]�?���?h[>*�?βH�C�/?'<z�8��JZ�hS�)	�=̻?T�?����\�y<�]�=�'��MZ�=Δ�U�"��pǽ��6<�_\�[��=�8=>�����B�=5�9�� ��1�&��=�t�@�����;'/L�g�=�����3y=H��=��L��L       split_indices[$l#L       /                                                                                                                                                                        L       
split_type[$U#L       /                                               L       sum_hessian[$d#L       /C̀CÂ?A��3A�C�d�@��Aq�X@k�V@�pS?�mpC��e?��@ZY6@�;�A�u@&��?���?���@9��C�5A�?�GI@5�@d��@O��@j��@�	?���?�)bC��j?��(@
h�@���?�?H?��!@<w?�
�?��a@`��BבC��w?��?�K�@��S?�Ja?�9:@ DL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       47L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       ������ݾ�3)��p>{��:����
�� >.� �0����#[;*�2��o>��7��r��<;F=��:�L>���=�j ��1�=��ھ�1D>B�N�bn�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L                    L       idI �L       left_children[$l#L             ����   ����      	         ����      ��������      ��������������������������������L       loss_changes[$d#L       >Ι>7��    >+��    >��>2.�>B��>~�>"�    >�&�>ݬ,        >�Q>y��                                L       parents[$l#L       ���                                               	   	                        L       right_children[$l#L             ����   ����      
         ����      ��������      ��������������������������������L       split_conditions[$d#L       ?��?�*F��=e?p]�=��?T>���?-M�>�u[>��v�ΐ�?'��=��������q.?~�9��=�1�<�ͽ�Ձ<�D���nR=iw�����L       split_indices[$l#L                                                                                                     L       
split_type[$U#L                                L       sum_hessian[$d#L       C��tC�lT?��C�r�?�`C�pA Z�Cݖ�@l��AR?�E�C�"�A�?�Vx?�/@W |@�#�C�p%?�k�@z��@��?ѤB?�\�@h�?��|L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       25L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       #:���u^>M;l��#�b��Y�>���U�2>T���9�qDh>����oL>�:Խ���<�90���=g�>�m�6Is>eϽo:;�� �<uOP>tb���qL=61�=�þ4۽���>��νBR>�y��>����bh<L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       #                  L       idI �L       left_children[$l#L       #               	                  ����������������      ������������������������            !��������������������������������L       loss_changes[$d#L       #>8�>#a�>�b�>?H�=a�>�zD>��>?}�<��=�p=��                >��>��t                        >��>R�0>��z>�=n                                L       parents[$l#L       #���                                                           	   	   
   
                                    L       right_children[$l#L       #               
                  ����������������      ������������������������             "��������������������������������L       split_conditions[$d#L       #@*It?�����L.?�����]�aǦ>86|�d�<�kP?�q��"*�=�|
����>#L��া��?�9<�x=�O��Z��=z,���W��'|����+�?;>*?�t<#$��X�����=����i/~��ڼ=��̻��$L       split_indices[$l#L       #                                                                                                                              L       
split_type[$U#L       #                                   L       sum_hessian[$d#L       #C7'�C1i@���C+�8@��/@)��@YsQC(��@S��@ܢ@6/�?� �?�*�@
��?��2B��B���?��?�n?�A�?�wg?��e?��B�@��uBX�zA���B�\�@�T%?��@P
dB9*�@��~@���A�sL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       35L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       :t���h;Y�1�H@���V�>�9:Ť~���<a�=�Q�� 5�w�v;�9��j^������c��Q�-��Q�<@T=&��m��?��;��J>Z�־Z����=i-����<�		L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L                      L       idI �L       left_children[$l#L                      	����      ������������      ����������������            ����   ������������������������L       loss_changes[$d#L       >��=&w�>=(B=�)�=�d    >���<�1�            =�*�>.��                ?j�?XS�?Kcb>�:�    >Y��                        L       parents[$l#L       ���                                                                                      L       right_children[$l#L                      
����      ������������      ����������������            ����   ������������������������L       split_conditions[$d#L       ��n���ʾց�?Pw��d�=�@���8\���k;�d�=ʒ�: @>�ڿOzo���,�ʿ���Dʻ{�j�[��M��?y�6?n��>)�O?�C�=�NN��Y߽��<2л�&&<�L       split_indices[$l#L                                                                                                              L       
split_type[$U#L                                    L       sum_hessian[$d#L       C���@��dC��L@`�@%?�ߥC�m@�
?��2?�Z�?��@O/C�q?�Ƨ?��l@ �7?�ӾA�-�C�.1A�fA(B�?�C�B�A��@�A�@��C@IC)TCCG0�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       29L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       )�αv:}�2���8=�����پ+\�=����A�n>Q-��p��;����o����>��S��Wf>�sy����>s�{��wi�G�=U�'>φ)��1x��4��t�>����������?:� �;��o��U�>D��1d>�>�1�>��=���;�v=���=zd`��kaL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       )                     L       idI �L       left_children[$l#L       )               	   ��������            ����   ��������                  !������������   #����   %   '������������������������������������������������L       loss_changes[$d#L       )>T�=�z�>�>�/[>� R=��H        >�l�?)7�>��F=�8    >�gT        =N� >F6>>��C=���>Z�:�4             =ZL`    >5!�>_�                                                L       parents[$l#L       )���                                               	   	   
   
                                                                  L       right_children[$l#L       )               
   ��������            ����   ��������                   "������������   $����   &   (������������������������������������������������L       split_conditions[$d#L       )?
ڿ�J&>����)��y>��V�<݃)�h�>�L@�����i�U<�0꽹�>�/����=�$+�U�?�tN�f���9��rI������������E�;�l��"K�[��[��:�
��3�=k׈�.;E=5J�>�7=���<��:�Z��!i<�<:�;L       split_indices[$l#L       )                                                                                                                                                   L       
split_type[$U#L       )                                         L       sum_hessian[$d#L       )C�RYCߛ�A�EA�C�[�@�3?�9W?��<@�
@@���Cؘ@�3@ �=@���?��<?�w%@���@���C�:@(�T@5��@�c:?���@4��?�F%@l"�?�ɿ@�C�0(?�#Q?��W?Ӿ?�G�?���@1_�@|v?�LO?���?�V;BQ�C���L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       41L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       9:��u��?�=䑺����>�'�<�-{�Q��=�־}��=w�b<�>�>����O�:<�I��vGB�ރ�>�M�: ��<�����=�<˾\tS;ߡǾ��p>��<'�e��M=߫j�,N��6�>�'� '��E�<�R�+�[>Lo����Q�>CTu�"�@��|<�� �uܿ.!>*�K���~��5-> ��=�hi��ǲ=�x�>�X���;�P>m	�<�^L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       9                             L       idI �L       left_children[$l#L       9               	                  ��������                  !   #   %   '����������������   )   +   -��������������������   /������������   1   3����   5   7��������������������������������������������������������L       loss_changes[$d#L       9>F>I+�>�ͺ>(z0>�0�=���>(۳?	*�?D>�;6>H�%        =��>�GA>�5�> �>}�\>�>5�I=3��>?�%                >��?��>÷Z                    >���            =؊�>E-    <y�0>E�j                                                        L       parents[$l#L       9���                                                           	   	   
   
                                                                           "   "   &   &   '   '   )   )   *   *L       right_children[$l#L       9               
                  ��������                   "   $   &   (����������������   *   ,   .��������������������   0������������   2   4����   6   8��������������������������������������������������������L       split_conditions[$d#L       9>v�P���?� ����?�9?��V�k����4��hw^���@-�;�~�=˙s����6��k�R���A���8	>���@L�@ {޽�E�;-޽�C�=��˿�>u�+}"�0�����%>�~�@.�Թ޿�8�Mա=uS3�s�<�[F@	bd�CTM� ߧ�	1>�<�վ'(=L�'�������j=@�<��~���<��G>
으�Z����W=�9;.�L       split_indices[$l#L       9                                                                                                                                                                                                                 L       
split_type[$U#L       9                                                         L       sum_hessian[$d#L       9C5cqB� B�?�B�Q�A��@���Bq�HB�eBpA ڵAτ?���@>�f@ͮBi,mB=�@v�@�_nB^b@Sh@�(�@�-�?���?�L�?�Nu@33vB]�6A��:Am�e?�DJ?���@UU?�Q@
�BU�"?Ů�?��6@��a@F�@�
?��/@ɩBT��A�|	?�#
AU��?�s-B%��A@��?�4?��@���?���?�@p?�R�@OuBG��L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       57L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       /9��+�t};6ly�P�T=���m��<�<O����<�s��ζ~�T��>��<�_��0���O�LZ�>������>A�V>���>��;��u>6������;��h��~�=��>�8Ƽ��(<�d�?�">�0i<�Ǟ�
o��[�=A���8mz�Ǎ������=0���E㼋D�=ϱ�>���W�>+AtL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       /                        L       idI �L       left_children[$l#L       /            ����   	      ����            ��������   ����      ��������         !   #   %������������   '   )   +   -��������������������������������������������������������L       loss_changes[$d#L       />`�>e>+g�=��|    >��>�]�=K�    ?,@,?9N;���>��`        >���    >��=���        ?'�>��+?'��>��=T�`            >���?2�=<� >^J<                                                        L       parents[$l#L       /���                                               	   	   
   
                                                                                      L       right_children[$l#L       /            ����   
      ����            ��������   ����      ��������          "   $   &������������   (   *   ,   .��������������������������������������������������������L       split_conditions[$d#L       /�M��?��>;�?���<�ά=��>UI�;��/=��v?R���&��?�վ�Te<�հƿ#v�>�>Z>#�R>��=/`?z��?�C��;��E���ɮ<7-@=�����0�[�?|�G����?ܭ��&߽�nE<hC��]P-�-�C�R���<T8� ����<�;�=�O��<Ϛ=M��L       split_indices[$l#L       /                                                                                                                                                                           L       
split_type[$U#L       /                                               L       sum_hessian[$d#L       /C���@�s[C��@��w?���Ch�C&��@T�?Ľ�C`m�A��@DJC#�??��N@�ZC^��?�4D@���@��?���?�Q�C��A?&�B!ïC6�@���?�`�?��P?�1�C�bA@@�h;@��2B	�O@�CB�2�B��?���@]kA���B�L�@`��A��?�Nx@x):@@�3@]1L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       47L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       5���:�#]����;�I\���輗�����:�:>
�;-�<.D����<>�!�}A����;��P�Sy�>Ѣ�<Y�Ǿ��<4ڽ>7ؾ��lJ^;7r=��8:�F�>�Й����>O�k��a;�Z��$>�����m=�>�oS>���-#�iԺ>�X־u�%;���=U��CT>楟��澿�< �=�����>:���6��L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       5                           L       idI �L       left_children[$l#L       5               	                     ������������      ����         !   #��������   %   '   )����   +   -   /������������   1   3��������������������������������������������������������������������L       loss_changes[$d#L       5=���=�OR=���>Fќ>#T�=��t<���>~��>�;�>�%?{M=y�8            >5"?z    ?��<���>���><>~        =��T>��,>�BJ    = ��>��x=�F�            >Tm�>��$                                                                    L       parents[$l#L       5���                                                           	   	   
   
                                                                                 "   "   #   #L       right_children[$l#L       5               
                     ������������      ����          "   $��������   &   (   *����   ,   .   0������������   2   4��������������������������������������������������������������������L       split_conditions[$d#L       5?�	?ܭ�>�� ?Φ?�i������e ?�2 ��1+<=��=�f�����=/�¼�������[O���=��7�(K|�V$��R ��H�������9@��?��y>�=���[�4����>�(�篠����=�k�>�06�2�]=���='�H�9���Lp=�4��N�:����3��3>
c`�>@H��O�;: �<�ﱽ���=_��[>_L       split_indices[$l#L       5                                                                                                                                                                                               L       
split_type[$U#L       5                                                     L       sum_hessian[$d#L       5C�KCߌ�@��C�C;A�� @���@%�\C�7gA!z�A�:A F@]�?�Zx?�s�?���C���@��O@�@���@�"�@���@��G@	O�?���@>NA?�C�~�?�=�@eK�@��@9� @>�r?�g�?���@C-�@�k^?��?���?��@�+�@�Sp@��xC�gN?��Z@�?��n@F��?�:@?�7�?��E?�\�@p�@�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       53L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       19x@5�Y0�=T.¼3���G�>��b<���<'۽�ײ>���=vd���]>$;;��>O:+��^V=Ё�= ��O>� ��3K�ofl;��>z�3=~i~�"�J><:�>���R�¼�W�>��8��z����n>�=9�x>6��=�G>x`:�D�I:=�a[�W�>�-0�B�=�݈����>I��>���<�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       1                         L       idI �L       left_children[$l#L       1            ����   	         ��������                           !   #����   %��������   '   )����   +   -   /������������������������������������������������������������������������L       loss_changes[$d#L       1>�>L��>QIJ>      =5��>L">&�>�m:        >���>m�R>v;�j�>��J>oy>�j=�1 =�2D=�?9    >.Z�        >�(l>�    =���>��=\��                                                                        L       parents[$l#L       1���                                                                                                                                                  L       right_children[$l#L       1            ����   
         ��������                            "   $����   &��������   (   *����   ,   .   0������������������������������������������������������������������������L       split_conditions[$d#L       1?\Kb?+߆����r2���^>��P?ԼL?g(@J=�Ob<�x?�f�@0�����	1>>�!@!r?J��?�@^?�<�>������ۿp��=���<���?� �=�2�=�{����?��>��P������Ӹ>Sg<^�=#u&�c��=���9>���q7=m��4i=�6:�i�=<�=
��_}=qҋ=�h�<�L       split_indices[$l#L       1                                                                                                                                                                               L       
split_type[$U#L       1                                                 L       sum_hessian[$d#L       1C3?�C�^BX�C[?́^@`�VBK.B�YA��@��?��^Aߘ
@��HB׊9@ٽAĽ�@�C`Aɂ+@0��@�@,�}?�DB��0?��O?�+A�s@BV@��@{��A�]�@a#�?�|�?��0?�q6?�x�?�@J?���?��FB��_A���@
�?�<�?�p`?�w�@��A���@��@N�?��tL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       49L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       -9ׂ��y;X���E�d=��>��:�Kھ��7��-�>����ü0z=7��|��=��z���:���:��A>=�b��b
�`e�6>"ú��|>_�I>�@!�I�=����i��>��߾��)=�ེ�3>�����\W:SK;�)>{�<�|,=�:ݾ��>���>��<�F}L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       -                       L       idI �L       left_children[$l#L       -               	����   ����   ��������                        ����������������      !����   #   %   '   )   +��������������������������������������������������������L       loss_changes[$d#L       ->��>D�>���=�M><g    >w�    >:��        >�D�?S�<�R�=+�?��>մ�?w��?K�                ?$*,>��&    >�{�?2�?!��?@�O>�-�                                                        L       parents[$l#L       -���                                                                                                                                      L       right_children[$l#L       -               
����   ����   ��������                        ����������������       "����   $   &   (   *   ,��������������������������������������������������������L       split_conditions[$d#L       -�Ytݽ��<�X �����>U^�=п�>��нةv>͙=�<8�"�����B�q%}>��P���?jQ�����P?*t��Bs��kp�Zs�=CQF>�IO��`g=��[���
�'S >��=���?T^��e<� A��Mq=�|ݽ�i9}�9:�t�=����M�<�yֽ�R=��Y=���;Ⱥ�L       split_indices[$l#L       -                                                                                                                                                                  L       
split_type[$U#L       -                                             L       sum_hessian[$d#L       -C�hAxlC��U@��$@&?i?�7>C�#?�@�#�?��T?��}C�G�B�m�@<6@)A���C��YB�a�A�.�?�Cc?�5
?���?�MA��@���?�%�C�3Bo�)A�Y@�}A, �A^8�@k�?��@e��?�q2C�~�B0l4A|��A�5�AF�@�!�@91dA �'@,=�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       45L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       #��*�;=�ͽ��s9�E5>�q˾���<(��;-�٪j��$���0>{���`�:5e�>���=�g�;�j8��F���(=��z>`Ѣ�
�;�ae>�7n��l����低���_>n���88>��5<�G-=�yE��&fL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       #                  L       idI �L       left_children[$l#L       #            ����   	      ����������������      ����                        !������������������������������������������������L       loss_changes[$d#L       #> Q6>�;>�h�>�.�    >9"�>XxA>g��                >�f>{7�    >��m>LÞ>�z[>�ޮ=-��=��=j�=�~\                                                L       parents[$l#L       #���                                                                                                        L       right_children[$l#L       #            ����   
      ����������������      ����                         "������������������������������������������������L       split_conditions[$d#L       #?�G�?������?��Q=�����w ���$?z���s�:|��'m=�%?_O?-M�=���<Zz/?Q|�?'潱Y����ƾ�F?�.?�/:�A�=�u��������JP�޳?=��輷�=��;���<�^S����L       split_indices[$l#L       #                                                                                                                                 L       
split_type[$U#L       #                                   L       sum_hessian[$d#L       #C�_C��A���C��?��@�ëA>/�C�g�?�9�?��~@A�?� �A��C�ZX@�@�@@���C̛\A���@R٢@T�@��@x&C���?��kAv��@���?�_@ �r?�"b?��[?�B�?���?�
~?���L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       35L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       C:�;����Y=
�,��0����=�$��˾�� �@>f;{h߾�yڽ��9=����R>�>7���3 #��>�,���<�8C=SƳ�t�-��1�>%/�<G�p�ug>����F����>�>r�"��;���=��8�r�>�[��`8>k醽��R=Չ�q�>��.=��l�>��\�hK*>�$i���=o�g>�n=+����C >��>��i���<�Y�$�b��[�=K��>�@d=��M�;�>rNb�՗=�1=EQt��f�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       C                                  L       idI �L       left_children[$l#L       C               	      ����                              !   #��������   %����   '   )   +   -����   /����   1   3   5��������������������   7����   9   ;   =   ?����   A������������������������������������������������������������������������������������L       loss_changes[$d#L       C=���>%Gc>�2>��>{��>#�z>�6    >G�>&��>3��>�.>o��>��>L�>l%>co�>2X=�D�        >^�    =�-�>�Ţ>�N�?m�    =,�    =�g�?��v?$�                    <�E-    >.ň<�@>S;~>���    >\Լ                                                                                    L       parents[$l#L       C���                                                     	   	   
   
                                                                                                           &   &   (   (   )   )   *   *   +   +   -   -L       right_children[$l#L       C               
      ����                               "   $��������   &����   (   *   ,   .����   0����   2   4   6��������������������   8����   :   <   >   @����   B������������������������������������������������������������������������������������L       split_conditions[$d#L       C�K�l�;*�>� ۿ���5 �oW2@R?��w��z��?s��@ª�3�r�XCe?,��@.�v�k~��2&->J�?�f ��|9<T����$���O�kLF����?2R?��x=�猾m�����g�ݾ�x�=�<��D��AP=��/��j�=���rk�= �a�=?H?�D?8L=�h�>�Gj=�+��1B<���>��<M����4>*�=�廙_�;�7��E�ݽ��#<tI�=�<��]�`j�=�b;�$3�=�C<l�%���L       split_indices[$l#L       C                                                                                                                                                                                                                                                 L       
split_type[$U#L       C                                                                   L       sum_hessian[$d#L       CC1qMB�߻B��BǾ�A)XA�3wB�?�8�BŲ@�US@��]@�Y�A���A��@q�l@�LiB�MG@Y�L@4�Y@H 	?��`@r(�?�c@��A���A���A��?�?@Ǭ?��B@/��A�B��v?��
@�?�h�?�"?���@K??��@j�LAR�A.�A��$?њ_A?�E
?���?���?�K#?��@@��?��@ma>B��l?��?��x?˒[@A�*?�#�A%�@'�AL�A�@?��F@ĥ�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       67L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       59��ӽ�q�;�	����>p�9�Qj=�㊾D��<�1�;��㾅�1�y�>�x3��q�Ӟ�>�����:��>�<�=�gl�۪�>�Ǿ$%D=_MF>Ϙ��7��
M�>��۾���=|�>��0�H�c>8(�;�c������5=�Yi>~���c���9&>��>ԫ;�&�<j۸���:���>yh��/弊�s�b��>����$�=�N�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       5                           L       idI �L       left_children[$l#L       5            ����   	                                    !����������������   #   %��������   '   )������������   +����   -����   /   1����   3��������������������������������������������������������L       loss_changes[$d#L       5=�=>���>If>���    >�4w>���>��>�c�>�b>��!?[5>Z =��?=^-=6��>`�<>��                >���>5x�        >��M>b��            >j��    >PB�    >'ݶ>���    =�K�                                                        L       parents[$l#L       5���                                                     	   	   
   
                                                                           !   !   #   #   $   $   &   &L       right_children[$l#L       5            ����   
                                     "����������������   $   &��������   (   *������������   ,����   .����   0   2����   4��������������������������������������������������������L       split_conditions[$d#L       5��n@\~?�p佁~~=��?��ؿzz?�O0?�N?ڈ?A�[�R��>]G>d?�}�C,@ p6?�mO=ԯ/<�₾��=쌉?��(@ ^=��� ��T���v��lv<��s=�Ծ���=\��?ӫ]��j�@I��L��=��*@��Ϊ�=-��=�3�G7�;��<���:O�=��о �#��j��=�#����g<�^�L       split_indices[$l#L       5                                                                                                                                                                                            L       
split_type[$U#L       5                                                     L       sum_hessian[$d#L       5C�SA �C�)A�7M?���C�nOAwV�AF�YA�@C�s�@}+�A
I@�c@ā)@��@>(@�2�C��;?��+?���@;�?���@��@]޲@VX@R��@6Ow@XET@9��?��@?�?@���?��C�)�?��@��U@<�S?�p�@�=?��>?���?�b�?�'�@7�Q@>-C��@!�@.�?¤?� U?�^R?�Y�?���L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       53L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       '�Af�:Y��,8x;��Y�\Fݻ�rԾjA7: 8�>��]��b~����;jD�c4����>���S�G<��:\@2>]}(��Is�L��>�u�$?�?q>I]�=?���q_=�����%�<���}e�>�X�u��<O>����>������3>�`hL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       '                    L       idI �L       left_children[$l#L       '               	��������         ����                        ��������������������   !   #����   %��������������������������������������������L       loss_changes[$d#L       '=�M=�E=$�?3�>���        >��>��>���    >m�=�8�=��=��0>�&�>�	�>��?
��                    >j[�>saq    ?H�                                            L       parents[$l#L       '���                                               	   	                                                                  L       right_children[$l#L       '               
��������         ����                         ��������������������   "   $����   &��������������������������������������������L       split_conditions[$d#L       '?��R?΄���r?��'k[��#e����?��?e�m?먟��1?��c���D+�?�۸�)
3=�h(�k>$v ���uo�=�Z�E3>6j�?�k~�1R��Tپ����`�;�L��	�=�6}��l��Ԯ�=��;J�=����>=���L       split_indices[$l#L       '                                                                                                                                             L       
split_type[$U#L       '                                       L       sum_hessian[$d#L       'CߎC��1@Jq�C�rMB7 ?���@�C�.J@� �B{�@+�C��@��@�@���@��\A�<fC��@���@H{!?���?�f�?�r&?�|�@3V�@DB�@Q�(A�SJ?ޑ�C"źCg�@:�;?��b?���?� �?�*?���A�QA�BL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       39L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       #:�3�;�}l�'=�9���>�y���"=���7�;=�С�_�L>�_/��)����>H��:�>[�����>߂����B��Jh>w�t;Kl��Ӑ>�h��G;�nA8=Tx�;���Y�>�ؽ�1j=N�.>�}�ɧ>8��L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       #                  L       idI �L       left_children[$l#L       #               	��������                        ����������������      ��������      !����������������������������������������L       loss_changes[$d#L       #=�[>�s>u>؆>:E!        >ϙn>}��>�Q�>��v>k�v>Lx�>���=І+                >�41>Z��        =�dh>=�                                        L       parents[$l#L       #���                                               	   	   
   
                                                L       right_children[$l#L       #               
��������                        ����������������      ��������       "����������������������������������������L       split_conditions[$d#L       #?:h�@��?�C?��ھRߞ���)<7B�?�ɾ?}�?���>86|?��z�o�쾁Ҹ�"=�=�ͭ���\>"���?J�>.�G:t�����B?��轎��<~�::��3��D�=����<x48=�c����=]��L       split_indices[$l#L       #                                                                                                                           L       
split_type[$U#L       #                                   L       sum_hessian[$d#L       #C.�C+�4@Cx�C&9�@�H�?�6�?ɻ C�&A�6?@ �@Fp�Cb�@��A��@r}4?�8�?�	N?��?��>C
��@3Y5?ԭ^@)��@�_sA�w@��?ǷRC�@���?⃜?�.�@m�@�(�@̫�@!L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       35L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       98��H=3�.��L�n�I>��Q�� ��y�^=YG}�g�q�
4�>�y1�qmX=�<c�Q?�P>s/澖�?#�>
�L��~���
>L(6;��M=��ս��Z���߻���>�&�s����;#���F<�J>��d��*S�3{�=cDt�G�F>5����[=��N��8�8�>l���k���P=�x>��9����>��g�P��94>hһq�%��>�Lt<�KtL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       9                             L       idI �L       left_children[$l#L       9               	����         ����            ��������   ����            !   #   %   '   )   +��������   -   /��������   1   3   5   7��������������������������������������������������������������������������������L       loss_changes[$d#L       9>i�?��>�Z+?5�?4{�    > �/?3�J>��    >���?/�>�4�>Ԁ�        >���    =�

>��.>͚�>�?m�?P$>��<=���>��2        ?��?@1        >K� >�?b >��6                                                                                L       parents[$l#L       9���                                                     
   
                                                                                             !   !   "   "   #   #   $   $L       right_children[$l#L       9               
����         ����            ��������   ����             "   $   &   (   *   ,��������   .   0��������   2   4   6   8��������������������������������������������������������������������������������L       split_conditions[$d#L       9�X�.�[�W���]mZ�NV���3�?^�4�^@D>?�%ض>��7?Q'z�W4��0��>#�=�銿[�D>C��?���-'��"vj?�<=��=Q�H?m�8�09�=���=������?�0�(�^�'ň<m�=����
��]�2?��սo�U=Y�Y��mM<�5����;w4=�����yt��S�=�=�䫻׸=�:|�.-��w�=)����-�2�4=���;�Z�L       split_indices[$l#L       9                                                                                                                                                                                                              L       
split_type[$U#L       9                                                         L       sum_hessian[$d#L       9C�y�B_ �C���B>ӖA5@i�C�w B�A/�"?�x�@��C�1SB��B��?�t#?��HAHy@{ѻ@F7C�#w@�v�A&_Bh��A�c�AK�N@�H�@(��?�7?�UjA��Cu�^@�?ߣ�@�@�@�� A:�pB9�2@��A���@�w@��@��+@=&�?��l?��A/�@���@��Cnu@�'.?�f??�X\@?��Aя@0_�@��B"*�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       57L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       =�M^�:�������;٨��V��<ܸ�S_":��>�L"�ذ`=�ļ>a{��f�=U���/;��R�^>����s�5>s��>�]����=��z�YL������N;K�>R�Ƚ�Q��&�>�/\> ��>c�˽/�>Ǵ�=�ѽ2p�>��\���p>>J�ѽ���;�밾"m
>����h[=�͛�i>Ll�=F��=�<�>��>�~F�W�|��RP���������W��9 >s<�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       =                               L       idI �L       left_children[$l#L       =               	                  ����   ����            ����   !   #   %   '   )������������   +   -   /��������   1   3����   5   7��������   9   ;��������������������������������������������������������������������������������L       loss_changes[$d#L       ==�&�=昆>&��?Qm>�^�>{>]��>sߴ>��>��>�m�    >�)    ;�c >L��=��\=_��    =���>��>��>�(=�?�            >	�f>�>��        ;�� :�     =�V
>���        <�t=d��                                                                                L       parents[$l#L       =���                                                           	   	   
   
                                                                                         !   !   #   #   $   $   '   '   (   (L       right_children[$l#L       =               
                  ����   ����             ����   "   $   &   (   *������������   ,   .   0��������   2   4����   6   8��������   :   <��������������������������������������������������������������������������������L       split_conditions[$d#L       =?� ?΄��>?� @5��?�H4�4?��L=�C�4@@�n=�I�=���<�`�����?�Ę>�ŵ�����c�@lʿP��'��@Q�??
X��9�����=+?��>k�]���<��.?>O�?���@�R��?��r�!�˼V �>�8���C�	>=s'b����:��m�B�@=�Ľ�i�=�����=uO_<nd&<��=���=�dT��M����a�ŉM��k����ϻ��'=��@L       split_indices[$l#L       =                                                                                                                                                                                                                          L       
split_type[$U#L       =                                                             L       sum_hessian[$d#L       =Cݬ�C�Z�A*3+C�V�B!@�6@�Y C�(Y@˘Aǵ(A�?�D3@z�S?�N�@c
�C���@���@���?��`@J��A�_@s�H@�f5@��?��?���@iC���@w�@9��?ƞ�@��@��@
0�?���@1�A���?��J@��@0��@ "�?��?�m�C��@�6�@2��?���?���?�ѳ?�8?��?�T�?�
?��?���@�d�AU??�n?��?�/?�5�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       61L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       1:�L:�7�=UM�޾g���!>n�5<�'�:�����=�N$>�n��L>-T��> �m�q�%<��<�F�s�>��O��u<8섽�ӻ�<V3>y�W�}�����>5�T��7��>vf>�r�2�t����>ׅ�=NF�!��>	�;�M>ro��?�=� �>�7ǽE
a=e��O1"��C�>�:=�]�>�*�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       1                         L       idI �L       left_children[$l#L       1            ����   	         ��������                           !   #   %   '����   )������������   +   -   /������������������������������������������������������������������������L       loss_changes[$d#L       1=��>�1>!��=��&    <�K >B�>M�b>��        >dNr>Bt�>+��>�1�<�0�>>n&=��L=���=�><>�    >Ku*            =S�6>N�H;���                                                                        L       parents[$l#L       1���                                                                                                                                                  L       right_children[$l#L       1            ����   
         ��������                            "   $   &   (����   *������������   ,   .   0������������������������������������������������������������������������L       split_conditions[$d#L       1?G�?+߆��>��h����?��|?ԼL>��i?'�<���=��Q?�ݤ@0����n=�޿>��?�@�?aP�?�@^?�<�@ �?��9?���b?�h������Y=Y����L?��?�@^�V���֎e>P(<wI!�Bx=$|�:�)8=�uμ�Lw<�41=�܉�lr�<9G+�x�]��`=-��<�=�=�̟L       split_indices[$l#L       1                                                                                                                                                                              L       
split_type[$U#L       1                                                 L       sum_hessian[$d#L       1C-�C
�,B��C	GD?�s�@P��A�*C6�A�?���?�cA���@�E�B��T@�۵@}�c@�RjA�r�@$i�@-L@!]�B���A��?���@��w?��@-|?�=@"�A�`�@8�p?�
�?��-?���?�p�?�d%?�W�B��,?�/WA�@K�L@�@T?���?��L?��A|�@���?��?؁�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       49L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       7���u��;)	�K+=�GU�	�N=B����;�l^��վ��g=�-޽<r��j
f���ƽ�� :�_b>s2��7оi9S=z�O��Z��N���<��;�!p>��V=Q���ɺ>�}a����il�>�Đ��U ��y�<8��d�q��Y˽�<� p�̎i>�����Q`=�?�>Ig���� �$>������W�Ү�b>�(�8T>�����|>m�=L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       7                            L       idI �L       left_children[$l#L       7            ����   	      ����   ����      ��������                  ����   !   #   %   '   )   +   -   /   1   3   5����������������������������������������������������������������������������������������L       loss_changes[$d#L       7>�T=��t>I�=��J    >ϫP>s�<�F�    >o�    >��?	%�        >�{�>G�?:J�?8��>�b(>�l�    >bsd=�a�>G"�?"�>�4?��>��>�P>j�V>��W>��                                                                                        L       parents[$l#L       7���                                               	   	                                                                                                                    L       right_children[$l#L       7            ����   
      ����   ����      ��������                   ����   "   $   &   (   *   ,   .   0   2   4   6����������������������������������������������������������������������������������������L       split_conditions[$d#L       7�M��?��?0\�?���<�� ?.�?�
�4TT:��>�����|?��L����l���U��e��?\��@q�<��?C�X�nܽ�a�����M��P�V6�?)ν�g,?��ҿ={>?
X?*~V>ô��^�;]���>w��8��A;�Z!��w�>e���.t<ڳ=qW��/�¼@��=�@q��ݜ� �k���?="�0�"C�=���3k�=���L       split_indices[$l#L       7                                                                                                                                                                                                        L       
split_type[$U#L       7                                                       L       sum_hessian[$d#L       7C�k�@���C��@��?�baC�	�B�>?@A�?�EC�=�?���B��3A�42?���@t0AlF�C��eB ��Bg�AY:A��@��AH	"@�8�C���A"��A��;A��{@�~x@l-�@���@�{;A%Q�?�*�A.#�@��@ ŌB���C4ǖ@G]�@�@�4A�@��A���@
�@�4�?�s�@s�@5��@'�R?�0�@���A
�|?� xL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       55L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       ��5�:h���ST�:�s%�g��c;^(�>�I�6mg�=��P>��~��K�;f�ཡTt>����Wݾ�2�>~�����L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L                 L       idI �L       left_children[$l#L             ����   ��������      	      ����      ������������������������L       loss_changes[$d#L       =�,=���    =̪u        >�et<�`>�ڗ=�7    >E�>ψ�                        L       parents[$l#L       ���                                         	   	            L       right_children[$l#L             ����   ��������      
      ����      ������������������������L       split_conditions[$d#L       ?���@,�=�}�"�p������=��o�|��겿m����J=�˿��j������=�Y���6=��p=�q��袨L       split_indices[$l#L                                                                              L       
split_type[$U#L                          L       sum_hessian[$d#L       C��@C��?�V�Cڔ�?�+�@E�C�
�@��TC��@w'?��@�D0CԆ�?�2?��?Ԁ�@TG�@�h`Cѱ)L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       19L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       M;(/]��#�=r������
�=��,�A�=��Ӽ����(���]=Oi>���ƣ=<=y���>S���Z7�{��3> &[���<�<c=��@�am��=��b>��p;�S�Q�=��>��<��e���=�-�7%R>	�=��M�^2�>Y�����<��Y>��Խ�1T=�ʔ�������>�ˎ�|8����>z>��X]��c3��wh=�Y�>���<�Ђ>n�o�i!`��{���9�����?~>w_~���j=�W����>赾1K!>��i�#�e��H>����=�E�+��>"bl��H�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       M                                       L       idI �L       left_children[$l#L       M               	                     ����               !   #   %   '��������   )   +   -   /����   1   3   5   7   9   ;����   =   ?����������������   A����   C   E   G   I��������   K������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       M=�V>�u=���=�*�>=3�>�{=�?�>��n>�r�=�t>/F=��    >Ԡ>�(>Q�:>^ʆ>ћ�=�I�=շ=vz�        >� �>=�>h�>b:�    >�=���<v5�>;,t>��)<�@    >��c=�:�                >+5S    >).v>c��=��=�/�        >J��                                                                                                            L       parents[$l#L       M���                                                           	   	   
   
                                                                                                                 !   !   #   #   $   $   )   )   +   +   ,   ,   -   -   .   .   1   1L       right_children[$l#L       M               
                     ����                "   $   &   (��������   *   ,   .   0����   2   4   6   8   :   <����   >   @����������������   B����   D   F   H   J��������   L������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       M�%Ʉ�;*�>� ۿ{\�5 ?©&�&�1�`� �f�K?s��@ª�o��=��U?���>���Wy��}����:M�>J�?�f ���;�{��oF?-��?��2?���=���@R�nh���&>ܙ��#V�� =���v�Խ�.[<�ý�Q�=���=�A(�=�82��B�?����f<:m�=�Z��5�D=��=�&��=�����(�=5�>dz;�-i=����Ծ �ǽ>��9aj����=�l��;�<��w�r�=;@�T��=�j~�Dj༰���I<�S�ND�=B܂�½�L       split_indices[$l#L       M                                                                                                                                                                                                                                                                                    L       
split_type[$U#L       M                                                                             L       sum_hessian[$d#L       MC+�B�śB�CBĈ(A�A�5�B.QAM�;B��@���@o�tAف@-�oA\{�A��@��'@�|N@��
B�� @Oi@(�z@*UP?�HA���A sA#��@br?�Q�A�i�@%(�@J�W@M�@y��@R�_?�jB�Ʃ@��j?�T3@]O?��?�r$AP��@�T@��@8�@I��@�(�@ ѕ?�m�A��?��?��?���?��?��@?�?��$@�}?�x�?���?�*6B�ѯ?�>�@7��@!�A@�K?�+>@�=?�2�?���?�@i@��@:�@e�kA^n�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       77L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       Q�tLT=��&2|<�f�>ݦw�N��KbK=O�r��'=s��?$z*��=t=��དྷS�<J�O<br->j�>Aؾƥ`���5�	R8>�J&��^\>-���L>v���S��=B]��C�c�ł�>��*�a�>�)P>f�*���=�����T=i�f�gG?6������Hkؾ��Y?�=ٹD=�vh��t޻Nh�>�T%>�'4���5>�签�+���>ߢ�����=�C�>V<>�nQ���,�T��^S>��?�7>���=z�?�;��=���
�∹>o�;�,�]�=a�? �7����>�a�;ۣ�>�8��CK;��L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       Q                                         L       idI �L       left_children[$l#L       Q               	            ��������                        !   #��������   %   '   )   +   -   /   1   3   5   7   9����   ;   =����   ?����   A   C   E   G   I   K   M   O����������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       Q>�f?),?>�t�>��>��0>�;�>�Ѡ>�r?��Z        >�(N>n�2?�K?a�>��:>ȱ?Nba?U �>��        =�S�?��P?+O@?��>���?�8?w
�?)Z�>��>MV�;8W     <��@>���    >i>�    ? '�>?PK>р�?L4�>d��?eѮ?Z�?f�                                                                                                                                        L       parents[$l#L       Q���                                                                                                                                                                                     "   "   #   #   %   %   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .L       right_children[$l#L       Q               
            ��������                         "   $��������   &   (   *   ,   .   0   2   4   6   8   :����   <   >����   @����   B   D   F   H   J   L   N   P����������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       Q�R�s�Ss�L��?��6?���>�Ӭ����?Uh�9��<�J�>E_f>��c?�Z������X�.<Fx�UP��V6�Nj�$�=ǌ.?"�������9���0�!�˿[��)��?x~n�Y�?É0�[k�=�i�?��J?�@^�"�?@1½����������?�R��+?%���gȿ&�G���w�=���=�ȥ��Y=��i��'�:>.[���<<�2=��>ud�8>
�Ofe�8�=�M��fv=�Z�<�Q�>��O��|J������=R�:�h&�)�p<�Pt>@橽��N=�uP;Ȥ=�D�j	�;ţL       split_indices[$l#L       Q                                                                                                                                                                                                                                                                                                     L       
split_type[$U#L       Q                                                                                 L       sum_hessian[$d#L       QC���B�ΈC��B��P@AgAgw�C�OHBb>�AM|?�%7?���A �@��MB[_Cu��B?"A�~@���@�T*@���@>0�?ŴR@OrA��B5$�AlIxCg7B&��@�[@��@��@5�}@h"?��V@��@�m�?��@w
?��@�`@��B+�A��@|�DA-�B;C@��B,@���?�ԟ@�%�?��w?�^<?��@@��?�=9?�1�?��4@#�@~�?���@Q~�??��?��L?�{?��F@�l?�AAԇVA��@��@��?��W@7�@M�@�sA���@�)A�V{C&�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       81L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       ?�C ;>4n���(���<Q�����=��&�Y�M��1�=�t6;n��=���Cd�>�#޽ՠ����><׽pYտ$p�>^z�I���y|q;�>P����3�� ����= �ڽ�W�jL>�ٺ�M>��(����>>�K��GR<n>���;JI���������M�->����F��eY�>b$M��	�e��?�c�tiH=O[�>�2߾1C��6�ξ�
�>���_C����>�·����<��>_͞��EL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       ?                                L       idI �L       left_children[$l#L       ?               	                        ��������      ��������      !   #   %������������   '   )   +   -   /   1   3   5   7��������   9   ;   =��������������������������������������������������������������������������������������������L       loss_changes[$d#L       ?=�Z�>�>2s`?,�>��>U�Z>a��>���>��>��>��P=��s> �        >��?�e�        ?�4?QF�>C��>��            >�]?|�?E8?OO?T�V=��F>��>.&|>�        >h�@?��>�5                                                                                            L       parents[$l#L       ?���                                                           	   	   
   
                                                                                               !   !   "   "   %   %   &   &   '   'L       right_children[$l#L       ?               
                        ��������      ��������       "   $   &������������   (   *   ,   .   0   2   4   6   8��������   :   <   >��������������������������������������������������������������������������������������������L       split_conditions[$d#L       ?>]R�R�s>���Ss�G��Yq`>��?��6?���?�+-�Ep�ۃ�;=>d=�ĥ� -;�{��9�ȼ�5�ET�VWU?�!���ϿP�=zG�
��Zx��n���{��M�տUP��V6��D@�Č�?�9>��Y����;/F�y>,�EG@�	T����мw
�=�
q�]����#=��b���?��ˍ>'�D����<x�K=�	ٽT���[N��l�=�{���f�*�=�驽�&;.�=�H,���L       split_indices[$l#L       ?                                                                                                                                                                                                                                    L       
split_type[$U#L       ?                                                               L       sum_hessian[$d#L       ?CڙC��Aw@GB���C�q�AM��@&JB��@A�	A҅�C�IE@6IJA p?�|�?�eB�2AM/W?�?���A`_mAD�x@YQ�C���?��?���@��@�<vB$��BT�@��-@�f�@*7�A5�o@���@�0?���?�ݐ@MC��w@���@S'B&�A
,Y@�`�B��@5��@hr?��@���?ϳ�?��EA#�{?���@�@0�d@�;H@��?�&@�G@~��C���?���@��oL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       63L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       ;9�&Q�kN�=&:R��;��|y�>}�<=�
;�1A��z��ߞ�6n�=a� >Ҥ���P�=�C5�?�O>Р��X�=��轰�b>T�n= ��E��>~��4��:��4����>�Sz�Y�=�	���t��В>s�=����K�C=��-���>l��F���q>�@��V:��e=�6G>���=J��h�+�h�	>6�g>�6�����@A>/��>%��'E��`>��b�Aa�>j��L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       ;                              L       idI �L       left_children[$l#L       ;               	            ��������   ����                  ��������   !   #   %����   '   )   +   -��������   /   1   3��������   5   7   9��������������������������������������������������������������������������������L       loss_changes[$d#L       ;=�5g>H��>��>D\�=h>�>�}>o�V?�        =�}!    >��x>h�h>�}>�ñ>�q�>*�\        >#��>7��>2��    >�	=ľt=��>)�        >NBn>H% >�CQ        >��>G�.>���                                                                                L       parents[$l#L       ;���                                                                                                                                                             !   !   $   $   %   %   &   &L       right_children[$l#L       ;               
            ��������   ����                   ��������   "   $   &����   (   *   ,   .��������   0   2   4��������   6   8   :��������������������������������������������������������������������������������L       split_conditions[$d#L       ;?��?{S?:��?�j?'"��j\?�F�?-�?�0��?��Z�p?.�>=��m?oh>���>PXh�N���OX>��ټ�WC==�@-Z.���@o��X�l>�����?��|?U�v=�l��F@ª@,�?��4�to�<�+?��Q?�-�@8	��w=�G纻����F	<��> Y(<so}���罋��=[�=�u��������=S1l=n�����,��=�ݽh�=�ċL       split_indices[$l#L       ;                                                                                                                                                                                                                        L       
split_type[$U#L       ;                                                           L       sum_hessian[$d#L       ;C)\B�P0B2�B�=m@"XK@�r�B ��B��DA2yK?���?���@.b�?�A՘�AV�B�
KAO�@��4@�#a?��%?�� A�}N@�m�A:�?���B���@d	x@�$kA	�?���@��@D�U@_nA�'�?�VZ?��@��@���@�3B��?�<Z?�:Y@#�L?�0�@F0]@��?��<?��?��?���?�3-@�a*A=?�&@���?���@�?7@-V?� L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       59L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       C:aC�G�;<�(ܾ��m� ��=����m������2z>�QJ�<�<� �>�\\��>	Uf�@�����\>!�潎l=���?
7�,��>ώ�g'>���>�婾�1�>nˠ�S)�>�k=�k&=���p,v�a��=g�F>����ǡ,�J/�>|o�>��n��2R�8�?K����y�_~�\�>��Ӿ_�V���ؾj>CC��ϡ�>��]���$=M�ݾ�轀�e>�F`���>�u���g����w=�>��L=���>�+/=u@^L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       C                                  L       idI �L       left_children[$l#L       C               	      ������������                           ��������   !   #   %   '   )   +   -   /����   1   3   5   7   9����   ;   =   ?   A������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       C>&>��R>��5=p>�Ȅ?���?u�            >���?)�^=애?��?Z�?p��>�	>��R?J�\        >��>с�? �>k/>�i>A?d�>�G�    ?��?6�d?a2�>�qt>��3    >�l�>sq�<��>A��                                                                                                            L       parents[$l#L       C���                                               
   
                                                                                                                       !   !   "   "   $   $   %   %   &   &   '   'L       right_children[$l#L       C               
      ������������                            ��������   "   $   &   (   *   ,   .   0����   2   4   6   8   :����   <   >   @   B������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       C>���g��!zT?�>x�e"y�&�þq%}��A+�U��>�-�^s�?if\>�ŵ?le?*t�L@��Z~��W�O�\�<܏^>%ۭ?7x�?��>�3?�^0�Nc�?R�h?c8�T��>�t�a2I�c��?��J����?�3�=޿�����>��?KhT?�E��o��#w�>3'��|�"r���=�����f�㆝��v�=jQ��(�=�5���<w)p��̱��í=�Tt���=�'2��ֽŦ�<0��=���<��@=�3�<�&�L       split_indices[$l#L       C                                                                                                                                                                                                                                                   L       
split_type[$U#L       C                                                                   L       sum_hessian[$d#L       CC�1C��B�9�@b%�C�bBc��B~��@!$�?��?��rC���BH��@�ϧB$JA���AϤCy�A�mcA��j?���@�uB��@�R�A�aAOp�@��@�3�@�6Cr
2@Mb�A��	Al3wA[q^A��@�B�@HE^@@_�@�}�@4:lA7��?���?��?��'@��?�) ?�@��q@�~�Cj�<@5c�Az)A\@ͮ�@�Q�@��!A��A5X@l�@�?��?�ۭ@�c@&�S?�ˡ?��7A�@2�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       67L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       ?�e׹<S���\�;��W>������:Ъa��u<6��>�4����!=���2>.)���=�h��ϊ�=u��F
�> �?��>��G����\���g��S>��]�#������>kR���J��H|=��R;�M�>����<���>_�I��+�?�=��<.�Ҿ|��T�;>�5>��Uq�?>#�>(~@�2��6=��(�1����>�ZI>��?<��>�A߾H\���hq>�+O�y��5qL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       ?                                L       idI �L       left_children[$l#L       ?               	               ����                     !   #������������������������   %   '����   )   +������������   -   /   1   3   5����   7   9   ;   =��������������������������������������������������������������������������������L       loss_changes[$d#L       ?=��-?j�?��H>[�!?R�?b$?1��?/�j>��h=}�     >G8�>t�0>ڇ>?��>�S�?S?jy >��                        ?M�?0��    ?!�T>O+            ?	�?/Ȇ?��>��>�;(    >�%`?P?w?Y�x>�F�                                                                                L       parents[$l#L       ?���                                                           	   	                                                                           !   !   "   "   #   #   $   $   %   %   '   '   (   (   )   )   *   *L       right_children[$l#L       ?               
               ����                      "   $������������������������   &   (����   *   ,������������   .   0   2   4   6����   8   :   <   >��������������������������������������������������������������������������������L       split_conditions[$d#L       ?�/�=�y��wܿa��?�0�.	�=��$��O^�w>�`���(��<�Ž��UW =����N�?�@^�%`¾[>�=;4<>'��=����7h���<a�?�I?K�^�>($�D6F>�)п�N6����4V�=혿5���"=����<�~d�>�q����?��>Ƚ>�:�����'�=�?�=6����>d+=J1�VY���f�<��0�U8��=�9%=�p>bp5=�覽po:��J"=� Ƽ�y��@"L       split_indices[$l#L       ?                                                                                                                                                                                                                                      L       
split_type[$U#L       ?                                                               L       sum_hessian[$d#L       ?C��C~��C14JCxȋ@�KMA{�C'l�A*�@Cn�@�)�?���@=�g@��A�ɍC]@Ҳ�@���B��C!�?Ǒ4@T�7?�t?�6�?�qA@��_@�zHAN��@$�[C�@��?��5@;��?�q�Bz2�A[0{BLtB��@�m�@0�@��0Ag�C5�A��?��@SeA���B1�?��A>��A�#bA�B~�~BsT@�@�?ٚ4@ �F@��x@�AEC��@�4C@�S�@���L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       63L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       !9�OM;I��U���M�>	��;G�o��T�g$t>����,=�Mv�`�A���>;`���c>˜�o�9��ƾ�F>�Ƚ���~��� =�FM�-Iл�!�>Oy:> ���e�+>p�K<-nb�\�=�y�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       !                 L       idI �L       left_children[$l#L       !      ����         	                     ����������������            ������������������������������������������������L       loss_changes[$d#L       !=̜�=��Z    =��>2 > �=,�~>H1�>B�>,R�>3�5<yp=��                >4�|>_Jy>Pdd=�h                                                L       parents[$l#L       !���                                                     	   	   
   
                                    L       right_children[$l#L       !      ����         
                     ����������������             ������������������������������������������������L       split_conditions[$d#L       !?�VF@*It��C?����g�?���?�4D?��:>86|?Ԑ�? ��q!@�=`{A���D=�U鼏�5?�yȾ���'9;"=�������g=���O�-��(�=x��=@����M=�v�;P�� �<��kL       split_indices[$l#L       !                                                                                                                      L       
split_type[$U#L       !                                 L       sum_hessian[$d#L       !C&ۀC%��?�ԚC �D@��_CWu@���@�k@0�SC	��A�C@\�@�?��1?��?�2?�tC��@�]�Au��@T��?���?�L?�?�?�nVB���@K��?�0�@�Q\@���@��"@
]?�X�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       33L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       Y:�w��;_<�J;+%p��8t;,Zx>#(��E!q=.[��7.��F�=�����f�=�I|>����//����?��=d���(=Ӯ��sl=$i�<�>>Ȭ7�U�|=E�ܽ t�>pk�>��G�F}̽a�4>,w2�۪�>{̟��q�=]�_������н�K�>�ʾ�RI>o+=�u��r>��0<���A?�:�^���a����>#�8�h��=��V>�c��o�:�+<�z?��=�y��W��M�>Doؿ�O>��R<���=՟׾�p=���ӗ�w��>$g'>ͻ=���=�K�b�����R>�ٿ?4=�����̷>)�>Q>��a,��i��JL >nfE��k�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       Y                                             L       idI �L       left_children[$l#L       Y               	                                    !����   #   %   '   )   +   -   /   1   3   5   7��������   9   ;   =����   ?   A����������������   C����   E   G   I   K��������   M   O   Q   S   U   W����������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       Y>	z">x�>�*�>�N$>Ϧ�>��>�	<?�J?%��>�'h?��?A�]?H
�>v��>v+ ?2��?Ly"    ?���>��>�>��>7�>���>��`?T%$?	��>zD�>��i        ?#�T?K>Ҷ�    ?%��?���                >��8    >\e�>eTl>���?0�s        >�W?;H2?@>��q<��h>>Z�                                                                                                                                        L       parents[$l#L       Y���                                                           	   	   
   
                                                                                                                       !   !   #   #   $   $   )   )   +   +   ,   ,   -   -   .   .   1   1   2   2   3   3   4   4   5   5   6   6L       right_children[$l#L       Y               
                                     "����   $   &   (   *   ,   .   0   2   4   6   8��������   :   <   >����   @   B����������������   D����   F   H   J   L��������   N   P   R   T   V   X����������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       Y>��>	�p�*A+��\پVJ<�!�~>��J�ӂ!����?�aQ>p˚�&�þ�9�?H�?�����?}$�>'�3���>��h?z��?m�$?ԼL?if\�^���%`�?R4?^�>�8�>t��n0�?�~��f?���=�`>͙����`�����`�=���)xL=#��?��@5A¿W�O�\����>�����?tR?�?�1�u\�?�Q�=��ۨ��_�;���>=H�<�̾1m���U=k�j���>	d2<NB= ,��Ҫ=���[����=EH�=��k<�]�<�'㽈+����0=,�ҾK�=�h����=J�}={B��t���K��r��=�
*��NL       split_indices[$l#L       Y                                                                                                                                                                                                                                                                                                                             L       
split_type[$U#L       Y                                                                                         L       sum_hessian[$d#L       YC�1C�n�B�yECVgvB1�#B�e�A�N�B��3B�;�AzqB:�BO�wB8�AWJ@�2B�-�A+,�?�<�B�6�@��i@@�A	�A�pB;�@��+A�v-A�]	A��@��@�4I?�3�B��]A���A;�?��&@���B��V@���?��?�4�?�M*@��?���A�9[@��A�I�Aعl?�_�@uN�A<�A%�fA"cAA|V�@?��@�B�@6$�?��!A�fB+��?���AuH�@��@ck?��T@��@�B�*�?�	@�U�A�-q@h_P@Sܜ?���@;YA���AcAN\�@G0�@��AF�?�D�@�?�@]�AkA�?���?�.�?���@8�@U�uL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       89L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       A����<=Ƽ�F;���>�����#�|�<7ȍ����R�=�5?>5>侜�J=Q%���lA�r�^>�`��T��Ȏ�>Ll��*v=�c����<ǁa>�����;-=
;Ɛ�����-�=�g�<:0����y<>��>�}�+���&�����=��L��>���=��5��VȿA����=����5b>��=����������5��}�>d�p>��~���>�1���(�>�d'�QS�r�����/=H^�����L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       A                                 L       idI �L       left_children[$l#L       A            ����   	               ����            ����         !   #����   %   '   )   +   -   /   1   3   5��������   7   9   ;   =   ?������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       A=գq>�a�? ?�>�w�    >��>�Ȓ>l�w>�?A�)?0��    >�A�?c�Q?r	>Dӈ    >�~>�
x??|l?)c�    =̛�>� P=�m�>�Y>�._?8�>���>�?1�
        >�B?-�t>��(>�Ձ>6�                                                                                                            L       parents[$l#L       A���                                                     	   	   
   
                                                                                                         !   !   "   "   #   #   $   $   %   %L       right_children[$l#L       A            ����   
               ����            ����          "   $����   &   (   *   ,   .   0   2   4   6��������   8   :   <   >   @������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       A>��@Q�?�]�@�"=�8i�!�~=;���>AA�&�þ�9�=Y~���~x���#D�1�=�sV?if\�^���%`�?R4=;���FW����>Q7�'S����q�@���	l�W�O�\�;EԾj����?tR?���h=�+��a�<;K�u�C>zQ=����h$�4N���X<!s��sC=�AK<�)����9��B��D@��0�=�4�=��1�,S�>�V�~�=�ޖ�)�ʻ��ʽ�69<pq���/UL       split_indices[$l#L       A                                                                                                                                                                                                                                          L       
split_type[$U#L       A                                                                 L       sum_hessian[$d#L       AC��C��eB���C���?�vFBĂ�A*X�C�^/A(�BO̼B98�?�%~AS�B�Z�CO�A��?��B:�@��1A��2A��?��[Ab~B�+>@���@t��CK;@q@�ƛA�Q A،L?�j�@u+AD�A)�iA#��Ax#M@^��@��8B�'@�C�@���?��?��@*Bw��CYP?���?��?�Z!@��@;GA��=Ac#EAM�R@GW�@��AH,?���@�27@Xj�@��~A��?�ae?͡�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       65L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       9:�����==^=�j\��b>d�L<�.����>����z;�E<��>�`��9�<�!s=� +��O
=J��>�H�;����Ze�>+�Ƽ�:�>�QE< ,
�0x�>���>�X	�'��9�T>e&ؾ��g=Ӡ�y�a>�3��I�t<wΪ�W�8<����
�X�c���>�E��V۽�>��Ͻ�=�=EA�>ߏF�ì�ktu=�V�[����e=��C���(L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       9                             L       idI �L       left_children[$l#L       9               	                  ������������      ��������            !   #����   %����������������   '   )   +   -����   /   1   3   5   7������������������������������������������������������������������������L       loss_changes[$d#L       9=žg>�p>6��>�n|>���=??�> �n>Q�^<��@>���>���            >���>�@        >XS�?)�)?�5>�Z�>���    >Z��                >C��?-�
>BȈ>gW�    >�2�>�E>�ew=	4`>.�F                                                                        L       parents[$l#L       9���                                                           	   	   
   
                                                                             "   "   #   #   $   $   %   %   &   &L       right_children[$l#L       9               
                  ������������      ��������             "   $����   &����������������   (   *   ,   .����   0   2   4   6   8������������������������������������������������������������������������L       split_conditions[$d#L       9>v�P��'\?� �g�`�$Ŀ�V�k���nS��Q�����m;��=�j�_��6��oH���s<sR��p"���~>�X��,M¾gP�=�� ����S�2=�%y=��ؼII�F����~>^�:?\e���ԾO�c�Y�@e�>��f?����0o�0�>	����n�/O�=�K_��}Q<l�w>"ľ'����E�<0;���t߽���6vz<��꼵�L       split_indices[$l#L       9                                                                                                                                                                                                                  L       
split_type[$U#L       9                                                         L       sum_hessian[$d#L       9C%V�B��.Ban*A{sBǦ�@hRBR�@��E@�`�A��+B�m5?�!K@!��@ BJ�@�a@ L)?�I�@t�~Ad|wAeO�@�n�B~L�@7�BA�?��?���@'�!?�T�@�}w@�{vA.��@YO�?�� @��A(�B\�j@C)B5��@ɲ@���@%��@wiA
n�@5�?��9@v@i�Q@<n'?��-@�ԲBMN/@sC�?鬓?��oB��A4
%L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       57L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       [:����-<�H�<
�6��G�Y�=l�a>+�L�f�}�,�>�꽾��<z��4(=�U�>��f�b
���<KDu�mwݻ�e�>�X�G��=�����OG>*鄾O�{>ˬ�=�p��,X�?BbF>�M�W&$=G�����>j޼�|��=P��-=믴���W=<��R"�>�=��۾k�����<�J.=�E?	��~x>Ȗ<����o�>;�X��K��W=�Ɗ�?��>D'��� ];ܳ��[�H����Y<���=8����2>� <H�2>d�w�ٍ���C�>c�y<���>.>��C�'숾��->?�n>&�㾾�������>�	}� �v��>�t�?��=���L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       [                                              L       idI �L       left_children[$l#L       [               	               ����                     !   #   %   '����   )   +   -����   /   1   3������������   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U��������   W   Y��������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       [> �>��>���>�<[>��>ֵG?$��?���>W@�>���    ?q�x>��m>���?,c�??h�>7�U?&
@>�d"?fvT?��    ?^^]>�X>��    >��T>��<?d1            =�ɖ?��?^�i?�5?�g>��>}��>5��>���?P >�I�>s��?T�~>�^?1�o>p��>�        ?
w?8�                                                                                                                                                        L       parents[$l#L       [���                                                           	   	                                                                                                           !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   3   3   4   4L       right_children[$l#L       [               
               ����                      "   $   &   (����   *   ,   .����   0   2   4������������   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V��������   X   Z��������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       [������5�>]G��;?��?�%�H�徠���#v�>�2�=���f�<�5��l�{�@N��$8(��&� KZ���>�Ӭ��e >#����=���29�=M9?R���F<��/�Nе>iB�==Pþ��F@+�@CP�*tP��>?O��W� >�Y~?95�<!;��*�f��>΁+�Z�ھap��Wr�?�g�<+�>$���*��;��t���=a����;�(�=݆�f�=kb�� 8;kr�$;��qF�φ�;���<CԾ @�=�';p�==�LH��b��Q;=���;6���}�=�ӄ�I�=��]=f�=G�D��ϟ�
�@��C�=����A��9��=�%�>0$0=.dL       split_indices[$l#L       [                                                                                                                                                                                                                                                                                                                                      L       
split_type[$U#L       [                                                                                           L       sum_hessian[$d#L       [C�NVC6��C;�$C>B��B��HB��Av�C�B
J�?�d�A�|�BM�AR��BŲ�@�Jl@���A�!�B��A��AU@ ?�4�A���B�A��?���A5	�@��B���?��@?�m@��A;
@�sA��B��
A��ADJ@U�sA�Ac6aA�A6BA�u@���A%_.@�S@��#?�G@j�BK_�B*?� x@DA
ps@BfN@��H@0��@gK�A� @g�wB���@�}?��|?��%A-�?��@��?��(A�?��,AIZ|@��V@f�1A%�F?��6A�Aa�?��@�s�@-D�@��@���@=�C?�R+@60B?��@:~I@-a�B1�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       91L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       +��N�;*�2�]O����>f�+��W���6k:�he�Sk6��>���J�R<������R>%�h���$�.:>�" =�<��L��@G>��G����96K��V!�>����6��?ì>�
�$V�>�@4;��i>�#�=��|�	��<OA>��b.�偠>��#�H˳>��9�4?߾�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       +                      L       idI �L       left_children[$l#L       +               	   ����      ����               ��������   ����   ����      !   #����������������   %����������������   '   )��������������������������������L       loss_changes[$d#L       +=�c>�e�>g՝>JX�>g<d>�r�    >?s=M!@    =��>��Q>���=��>��&        =�Ĩ    >T�    >6.<>�H�=�kS                >d�N                >��>{I:                                L       parents[$l#L       +���                                                     
   
                                                               !   !   "   "L       right_children[$l#L       +               
   ����      ����               ��������   ����   ����       "   $����������������   &����������������   (   *��������������������������������L       split_conditions[$d#L       +?΄?� �'k[?��۾o��?먟����?�Ę?�8)��-��Ͷ�)
3?�ۑ@G�=	����_�3F?��<*6�1R��V��Z�?�˜�/��z�=˥��[0�>��?�.�E5+=��r:�>{�?5�J��~;x����B��	�-=�"+�p�q=�/x�XL�����L       split_indices[$l#L       +                                                                                                                                                          L       
split_type[$U#L       +                                           L       sum_hessian[$d#L       +C��
C`B�OC��;@��IA�|�@n�C���@i+?���@�!@���A��C��@�3a@�?�K�@s��?�5@50W@5�@��A��C��?���@5�M?���?���@:.?��?�[�?�"T?��A.�GA5Cx�B���?��y?���@�g�@f�Aj,@ǈL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       43L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       5:׈f�U�2=+�,��Wo�vkv>u�}<gT<X�'��_����P�=}66>�L6�6�<�����=л���<�dֽ���>F<��;g��h>R�:�u<l��,�����E>#�PzG>F��>mS��_��>�E����ݽeT=�#;���>����=m7���ç>H�'>�<E<�@j�~f����þ4�><<>�L�Ay�>sӾE�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       5                           L       idI �L       left_children[$l#L       5               	            ��������   ����                  ����������������   !   #   %   '   )   +   -��������   /��������   1   3����������������������������������������������������������������L       loss_changes[$d#L       5=��>8jn>t��>H�~<���=��=� �>BI�>2a        =��v    <��><�	>��>z�M>�#�>&��                >��>C�x>>��>�^t>��Q>�"�=��         >�Qb        >I=F>zG�                                                                L       parents[$l#L       5���                                                                                                                                                       #   #   $   $L       right_children[$l#L       5               
            ��������   ����                   ����������������   "   $   &   (   *   ,   .��������   0��������   2   4����������������������������������������������������������������L       split_conditions[$d#L       5?��?{S?:��=�V�?'"��j\?H.P���^?��[���v�z��?.�>=�(A��v��[P�[���.>�r�{�*���=m�}�`�˽�6�?���?����"��C?#�/��@��=nGy=�ep?2R=������?o>���:�u=������<�T˽���=p��=�{�;ڳ��������X��=a�;e)�h+�=?WʽlhNL       split_indices[$l#L       5                                                                                                                                                                                                 L       
split_type[$U#L       5                                                     L       sum_hessian[$d#L       5C"��BB,5�B���@Yn@��GB��B�p\A��Y?�?�?�sQ@(�?�@�JBs�B��5A���AWp�A��?�Z�?��o?���?��@�.�B�B��=A?�@t�Ag��AC�~?�cx?�n@��.@J92?�IMA��3A=VB�a ?��A@��@���@(��?��@�]H@�A[�@#�@���@HfAdl�@��rA$BW?ȝ�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       53L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       7:���μ;vs��\�=#��<>3J�(���{ǽz�;�b�=���=�-W��&���;<�YZ���>K��Ee>s('�zn��.���.o�v2]?$#�<�#L����=���=�r�>���y@w>�¼��O>�����=�]���};e=(��<�>��G����������=�7��g&>�V��-�>`�u�+n=�������k�>Q�	��=��z��XL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       7                            L       idI �L       left_children[$l#L       7            ����   	   ��������                                 !   #   %   '����   )����   +   -������������   /����   1   3����   5������������������������������������������������������������������������L       loss_changes[$d#L       7>�=�'<>�=-�,    >in�>���        >k=?��>zfN>��P?�?H>�8�>X}�>"d�>���?�>zmR>�;7?�w    >�Us    >i�>J�             =���    >D1h>�    >j(�                                                                        L       parents[$l#L       7���                                         	   	   
   
                                                                                                   !   !   "   "   $   $L       right_children[$l#L       7            ����   
   ��������                                  "   $   &   (����   *����   ,   .������������   0����   2   4����   6������������������������������������������������������������������������L       split_conditions[$d#L       7�M��?���>L �?sB�<Dd]����׹ν�Ǽ�.����:��!?@1�>p˚������T=�I>w��
�̾�ͮ>���/DԾ���̹�>D����@L��)\?W$�2%]=�'���=) ���Z�=��'�9.	?���1c?��"�$q=�9���ڼڊ��Y<<�u�?H�=����=���:4=�����Ⱦ�=z䱽%q�<�&�����L       split_indices[$l#L       7                                                                                                                                                                                                           L       
split_type[$U#L       7                                                       L       sum_hessian[$d#L       7C��&@���C���@op�?�b�C���BSz�@��?���C�ìA�}@��B5b�C&�C`�@��`A�&@+4`@�%�AʋB0SC�A!!b?��[CS2@E[�@�5A7��@���?���?���@=�@*�@��@W!?�(eB	C]�@-�G@���@�� B�Y�B.�?��?��\@�v@���?�>�?�<V?�W�@���?��.?�G�A�xcAEKwL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       55L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       #�� :����J�PS">�DA��==�7:�i�+�r��'��)�>_��L���$�=���>M�x���s>!ţ��<�?�>��|:g������GX>��J�4S>�ĭ>3����2<��@���$>M�k�z;�?Ɠ=��L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       #                  L       idI �L       left_children[$l#L       #            ����   	         ����      ����      ��������      ��������   ����      !����������������������������������������L       loss_changes[$d#L       #=�l�>S��=�Kd>��    >��F>�J>g>�D    >=�J=9�X    ?*�?j�        >���>��        >!�    ?4��>+�d                                        L       parents[$l#L       #���                                                     
   
                                                L       right_children[$l#L       #            ����   
         ����      ����      ��������      ��������   ����       "����������������������������������������L       split_conditions[$d#L       #?_�?T�1�?;B=��N?�g�<p�z?{S���ƽ��7?�x��u�.>���>��=w]���>�
J���;�L�=��/�/���>�9C?8>�X�=�7=V�����;�����=v�N��#�>1T�<��>L       split_indices[$l#L       #                                                                                                                                 L       
split_type[$U#L       #                                   L       sum_hessian[$d#L       #C�:"CȘ�AT(�CǨ ?��AAϸ@���C�j�@�W�@14@�V@ N�?�)&C��Av1?��:@Agz@7��@^��?�-�?�o�C��c@�uADX@F�?��"?�^�?�<y@	zCY=�C��@�l@�D?�v%?�c(L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       35L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       =;������<��P�(.��p�s�sdH=��=la���X>"	t���<o���.c>Q�<�n=�2~����>b9K�.�߾fm߼�<˽��x>BoN���a���
>�wQ�6�>��C�=[��<���>�ȸ�q����(c���k>4F*�r�>7�>>����P�>ִ�=�O�=(*H���^>wO�<�Ⱥ>�^ <ٙ�����Lp���ɾ��>��=� ��Zƶ=�k���=�����w	�>��t�d>=��<L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       =                               L       idI �L       left_children[$l#L       =               	         ����                  ��������   ����      !   #   %��������   '����   )   +����   -��������   /����   1����   3������������   5   7   9   ;����������������������������������������������������������������L       loss_changes[$d#L       ==Ӊ>�l>�>Fsb>W�>��>$@<���    =��>��>v<ی@>�\>WW�        ==��    <_S�=�0�>��'>�4        =n��    >�&�>؟8    =�F�        =��    >�	e    =�            =�0>ca>�(>>#�                                                                L       parents[$l#L       =���                                                     	   	   
   
                                                                                 !   !   #   #   %   %   )   )   *   *   +   +   ,   ,L       right_children[$l#L       =               
         ����                  ��������   ����       "   $   &��������   (����   *   ,����   .��������   0����   2����   4������������   6   8   :   <����������������������������������������������������������������L       split_conditions[$d#L       =��8�w���:R�������ǿH�!�(f���^���/7�4]ݿG���W�̾pp���w�c6=��	鷿uܼQ��`}�@W��>�`޿I�'���ۼ��-Wz�[6K�rC��A>�;��m�U_���𽪖�@(�=XT3���=\��=�u{��ǎ> ��<���<lgA��"����߼=�<�q�����uSҼ00%��M=��M<�'8��D=����e��՟��9)=�����<��L       split_indices[$l#L       =                                                                                                                                                                                                                        L       
split_type[$U#L       =                                                             L       sum_hessian[$d#L       =C �$Bh^B�@@��wBR��A���B��@	�@R�T@�^B=� AtX�@4�@���B��?��?�"�@{�9?��@�&B3٭A2@@�r�?��l?�>@V�z?�%;A�W?B|��?�<@9�2?�f�?�cNB/��?��KA�@>@G4	?�c�@��?��|A=L@�:dA��BX?�?��Q?�}B&eG@K9@��?�Q?��3?�i�@��b@�*5@6�3@��@ �@�L�A��B�YL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       61L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       I:�s���<@~k�[f������3<�뽾RhR>��>E�۽񠻺�0��v>���<S��y��=���>����fؾ�I����>��ὴf��ϟ^<�N;��>�ՙ�4��<��输k�<<zz��j�>����.H��D=3��#'w?Ű���>N�R�%��>.�?Iq�����)��c=ſ>�
�����V>N7��=�?d=�侉��>QPC����ܐ=�.@����]r��?n����>9|ν�hh>��̾��o��GP��H�>G�x=�y�>Y���W�=L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       I                                     L       idI �L       left_children[$l#L       I               	         ����                     ����   ����   !   #   %   '������������   )   +   -   /   1����   3   5   7   9   ;������������   =   ?����   A   C   E   G��������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       I>
{]>��X>O{�>�B?�>���?hR�>GFL    ?l�,>�Lt>��>{�>�+>��#>2�p    >��    >F_�>�
�>�l]>��            >H2 >��>�
�> d�> ��    >c��>���=0y�>�*T>��            >���>
�I    =���?��>��h?��                                                                                                        L       parents[$l#L       I���                                                     	   	   
   
                                                                                                     !   !   "   "   #   #   $   $   (   (   )   )   +   +   ,   ,   -   -   .   .L       right_children[$l#L       I               
         ����                     ����    ����   "   $   &   (������������   *   ,   .   0   2����   4   6   8   :   <������������   >   @����   B   D   F   H��������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       I>�]9�U�*�H�'@=�D>G�пS��@>�?�R=�#�� g>�G���K	?k@�=�PH�6K�?��<�i����i����>��">F�?KN��l����%�<8/:��l�Dmx>�ٴ>g�����d?������<(g�>iޙ�0a"?���><��>$ m��8=x"c�WA4�P�O>?$�?����a%⽱\t>@X�&6���I5=wv�c��>*�z<գ��@@={-���o<�7������	��&��Պ=^�ż��=�*��Xݼ�����$=o�]<&�Q��p�=�����c�L       split_indices[$l#L       I                                                                                                                                                                                                                                                                     L       
split_type[$U#L       I                                                                         L       sum_hessian[$d#L       IC���B���C���A��B�N�A��'C|~�A�&�?�B�A(��B|h?A[6�@���@��Cu�0Abj�?�A�@g�A G�B\V@@/ORA/b�@I�R?۟L?܋�@��A4��Cj��A?9�@Ý?��u@��@,@��lB-GA<��?�1�?�l�?��}Ae�@l�@$j�@�O�@͙�C/��Bj��@��Aű?��0?��
@�B�?�?�L�?��S@V�M?�mA��AR��@�#�@���@�x?��|?�2�?��
@P�?�X`@$H�@v�B�'�B��
B4�A�&4L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       73L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       )��q\8���ԥ;L����k;��z �]D#:j7>M9Ƅ�(�=�|ͻ��P=p/�>��s�,�O>RH4=.�����P�8>�||��Pd;di�����<���>�\���P�&z�>_�����=�3��{>��Y�7�=�o�>p���.�>Mg�*y =N? ƴL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       )                     L       idI �L       left_children[$l#L       )               	��������                  ��������         ����         !   #����   %   '������������������������������������������������������������L       loss_changes[$d#L       )=���=�� <��>0t�=�܏        >	��=��>�O>Ix<?-�>��        >E4>7*}>'�}    >���>5�P>���>�?�    >&��>4�                                                            L       parents[$l#L       )���                                               	   	   
   
                                                                  L       right_children[$l#L       )               
��������                  ��������         ����          "   $����   &   (������������������������������������������������������������L       split_conditions[$d#L       )?��R?ܭ����?�C��-8M��Ś���|�Z+z?���?�?��\3�?b]l�@��<��=��$=�I��^��a���y:�ʌ
���)�=�:�;����K�>�06��H����ǽG�=�2��"�7<��q����=�j�\��= �=�s1�48`=v|��L�4<wL�>�L       split_indices[$l#L       )                                                                                                                                                    L       
split_type[$U#L       )                                         L       sum_hessian[$d#L       )C͇EC��@5��C��vA��Q?��9?�b�C�[@X�aA(X�@�o�A�I|C���?��^?�Fe@���@��@#?B@g�KA�W�@�ƑA�	�C��*@A@@6Q@(5@ؓ?��?�q�A#6-A)y�?���@���A�V@��"@��=C�-A?�ю?�Y?��?��qL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       41L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       1��6��� �>	I�<�K�׈���>�?�;�ͳ>+e����<���n����>Ɔ����X<���c�i>�mu;��.�)�M����>{E��kh;�$�>x=�>�=������>\o�Z��=�Ǧ��?+<׸4<��$>��=���+'�<ܴƽ˼������2;���S,۽.,>2��>
1L�6������=��L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       1                         L       idI �L       left_children[$l#L       1               	                  ����������������   ����               !   #   %��������������������   '����   )   +��������   -   /������������������������������������������������L       loss_changes[$d#L       1=�p_=��9>-~�>- '>'�H;�M>�> �>P�>59�>�XG                >%�&    <�� =�l>Lj�>Y=�oH>�8�>"$�                    >u�|    >D<�>i�"        >��>�?w                                                L       parents[$l#L       1���                                                           	   	   
   
                                                                       #   #   $   $L       right_children[$l#L       1               
                  ����������������   ����                "   $   &��������������������   (����   *   ,��������   .   0������������������������������������������������L       split_conditions[$d#L       1@*It�d���L.>���?�9�6�н���>�WZ�׮��JA?�t�󮅺�m=�;)�������s���P>��@UT�/��>������^�2��=���=�;<��e�/�=9;�?�(=��>��>݄:;�;�=�9H?�6�?�>�<lw��{F�����0#p:���}i�P�=V��=%�½[2c���=�L       split_indices[$l#L       1                                                                                                                                                                                L       
split_type[$U#L       1                                                 L       sum_hessian[$d#L       1C�~C�@���B��0B�O�@ P@'U�B�_�@�GRBD�SA��?���?�7?���?��/B��?�@Fӑ@I�AC�(B��@��cA���B��@��@ X�?���?�j`?��A*d�?��rA�IJA�I?Α	@�BA_7A �Bh#�A.��@�D0@��DA!@���AiQI@���A8��@�@��=@;L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       49L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       79F�`�m0Y;��!�+��=^�f>p��;�&��I�t>,��>(���7�,�4<�����ʽݙ$>�V*��ػ�ׇ?;��
��{=:��[;n�=տ;��㽦��>uv�*��;v�N>�=������>�U���xȽsoa=��D<4����S_����>SB>D�e���I����=��=��#>���80=�WH<��>�����o�@�>+�߾m�%>��%�s�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       7                            L       idI �L       left_children[$l#L       7               	����      ����                        ����   ����   !   #   %����   '����   )����   +������������   -��������   /   1   3   5����������������������������������������������������������������L       loss_changes[$d#L       7>�>�2M>&>`>�-    >3͢>!�(    >�"M>���=�z
=�C>5��>T~|>>x8>�,    >yń    <�L�>c�Y>��"    >}:�    >P�$    >�l            >��        >7
.>��>V�> �V                                                                L       parents[$l#L       7���                                               	   	   
   
                                                                                         #   #   $   $   %   %   &   &L       right_children[$l#L       7               
����      ����                        ����    ����   "   $   &����   (����   *����   ,������������   .��������   0   2   4   6����������������������������������������������������������������L       split_conditions[$d#L       7� 5D?^�9�!=�@-F�?���=�Sa��n�4l�=O=�JA?�S�>�|?�p�>d�3�ؿ(�?���Q&?˰l�����;�?���,v0��"?bp0=<�[>�G�:�'���P"<�8Ľ��b=�3�;�����<���?��X>�C�O<��5j =lLz���%��xL<-�3<��>	6a�]�=4_;,O�=��轷@�g�=NT?����=��Ƽ9WvL       split_indices[$l#L       7                                                                                                                                                                                                      L       
split_type[$U#L       7                                                       L       sum_hessian[$d#L       7C�.�B|�C�JA��A��?嶡C�9�A��?�)!A)V�@��@���C�ݵ@BA.@��@?0�?��!@�1@��@�C��dA=*@W��@-@�?��zAA?��i@���?�ƛ?՚�?��R@��?�y�?�oC�j�A���@xQ�@�+X?��
?��U@��0@HL�?ߺb@z �@t/?�VeC��g?�>�@��`AXr.?�R
@.��@�0�?��L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       55L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       �%�=�U��ͽ�_�>�퉾E��9밝>�S>������;��>Q�~�.6���E>�v"��1)9��)=��$�n�w���4>,�L�����y�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L                   L       idI �L       left_children[$l#L                ����      	   ����������������      ������������         ����������������L       loss_changes[$d#L       =�i%>��>S�:    ;G�=��6>�;J                >cJ2>��@            >+�>��.>��                L       parents[$l#L       ���                                                                    L       right_children[$l#L                ����      
   ����������������      ������������         ����������������L       split_conditions[$d#L       �o�|�p�e�m������겿V�r�j��= ;�=�A�� :�n��|���it5���=ƍý�:��c��f�¿b����w�=Oz½�D��L       split_indices[$l#L                                                                                               L       
split_type[$U#L                              L       sum_hessian[$d#L       C�7[@ν6C��f@7N�@f+�@��CŰ?�t�?��(@6�i?��@�#IC�7�?Ȭx@W�V@T��C��!Ax��C��@f�AS��?�H�C��L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       23L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       A�<F�^�Q=U��;Կ����>\�<������<�'� 1�=7(6>���<D��;n�=0�Ӿ�=�I�>��@<6EȾ=�����>H�׽��>-o�<]b�G?���Ǩ�#1	>�s>f����5��q�=���>�ˉ��%�>~�=�z�/��=���>�n�����>	(}����>1q��J��������=�r�>Θ]��������<B�|����=� a�Zs�>4��1�=[;u=�`�>��i<����p��>�iŽ��L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       A                                 L       idI �L       left_children[$l#L       A               	                  ������������         ����         !   #   %   '   )   +   -   /����   1   3   5��������   7��������   9����   ;����   =   ?����������������������������������������������������������������������������������������L       loss_changes[$d#L       A=�4�>>�U=�1=��c>Jd=�e�=��X>]r>��>�F>u            =�*8>�SL>CF0    >_��>z��>��<� =�9�>t��=�w>:��>B.�>z�    >U�D>˴�>Q,        >_�        =�%    ;�>�    >0�x>=�6                                                                                        L       parents[$l#L       A���                                                           	   	   
   
                                                                                                   "   "   %   %   '   '   )   )   *   *L       right_children[$l#L       A               
                  ������������         ����          "   $   &   (   *   ,   .   0����   2   4   6��������   8��������   :����   <����   >   @����������������������������������������������������������������������������������������L       split_conditions[$d#L       A?Gļ�r2���ڿW�`@5
�u8�>�>���[&�V�5>�l@!r=�$�;'0�`�A�b�P�z�Կ�&=�^��H�?�D?�ƿ"s���>��P?ԼL��[O;�l�o�=�#W�Wy�=}�@J9n=
�=��>��=�iE<�`R@=�<����N�����?�ݤ@0����=T���� �>fȽ���<���=��
���'��);i�����@=yԽ�<=">m��;�<��=m=�x;�?ҽ�Y!=��S���L       split_indices[$l#L       A                                                                                                                                                                                                                                          L       
split_type[$U#L       A                                                                 L       sum_hessian[$d#L       AC��B�h�A��B�A�>�@9�2A���A���B�w7A��@«�?���?��{?�l�A�%�AF,�@�ĳ?ێzB��AU��@�`t@a�@g��@���A�CW@��)@�l�@��_?�aR@_=�B�A9��?�P�?��T@���?���?��6@S?�E�@J�+?��A��@���@�0@%zG@L,h@��?�#�@\��?�w?�?ҎB���A(�$?�$-@��7@ �P?���?��-?�S#?�32Au��@�@J�?�U�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       65L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       -9�|��М;��I��>8OM�ҩ�<s��f�h=��Zg�}e5>\��;�Ā��Z��Y�>�^����C�޺�>Qv���\νQZ>�{<@�j
�;��̾�}6�$��4�#>x;��;>�C)��":�z�/Uc;�7�>��;���=�S�e�@>��ؾk�s�e:4�i+���7=��VL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       -                       L       idI �L       left_children[$l#L       -            ����   	                                    !������������������������   #����   %��������������������   '   )��������   +��������������������������������L       loss_changes[$d#L       ->�^>n�e=���>�-�    >��>R�k=��>�a9>2b�<�h=�<:>6�=n"�=���=�M�>n�.=/��                        >.D    =��                    >厷<�P        >*�                                L       parents[$l#L       -���                                                     	   	   
   
                                                                 !   !   $   $L       right_children[$l#L       -            ����   
                                     "������������������������   $����   &��������������������   (   *��������   ,��������������������������������L       split_conditions[$d#L       -�ǮO@�,����?�7t=]+���Wk��Ŝ?[��?����?>���R~����3�e�`?[�ܿEB?�S�� g={[�����{8�=�F�;�&y��l;��n���u>��&�Y+=2Ԑ:�xG=��2���l?ݙ�?:�;��=�F�?Jd�<3q�����=�Sj���y���S��樺$U<��L       split_indices[$l#L       -                                                                                                                                                                 L       
split_type[$U#L       -                                             L       sum_hessian[$d#L       -C��A�LQC��LA��Z@'�A��C���A+��A�@��6@4$l@pBuC�@�o6@/]C@h�@���@��?�dp?�L�?��?���?���?���C�mR@:K@�l�?�U!?�ee?��}@��?�N@�I@1B�?�z�?��C��?�,#@oC?�9s@-�R?�
?�ևC��B!L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       45L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       !�H|:��ξM�=�`	�?�����p�V�*��q�>�	u�
�;=�q=��>�Ϝ�Pf=�~�=�?�Qp��۟���<>#[�>�9:���X�@>~�>iM8��V���y>WՅ����9>?=K�o'L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       !                 L       idI �L       left_children[$l#L       !               	������������         ��������   ����         ����            ����������������������������������������L       loss_changes[$d#L       !=�o�=��g<�<>�">FHO            ;�Q@>M8<>�?        =İ    >�]N>n+�>���    >r�B>���?,�>�DE                                        L       parents[$l#L       !���                                         	   	   
   
                                                L       right_children[$l#L       !               
������������         ��������   ����         ����             ����������������������������������������L       split_conditions[$d#L       !?��R�o�|����p�e��#V��n��M�����겾otο`�=;s=���C=壼�ǿg�D�X��X�=�Kj�,'�g��c'潁�Z=���=��"�����_=���+�*o=e|���p�L       split_indices[$l#L       !                                                                                                                           L       
split_type[$U#L       !                                 L       sum_hessian[$d#L       !C���C�_u@1�o@�lC�9�?��?�Q%@5�_@]�An�C��M?�TE?��`@�?���A���C��Q@�>N?݅A�0�@6v\AU��C�)�@� �?�w"A@�K@�9X?��m?�KA=x�?���Aw�C��0L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       33L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       ':�CĻ�X�=����O�/�h�>g��@�<?�E�r�=��~>�R�����>;h{�"k =��=���C��b8>��L�R.r�gH>�l>>���{^��X"=��s=�?�@�#<�=�*�A>�nw��H}>��o��R򾴸�>
�U=��<�>4�`�X�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       '                    L       idI �L       left_children[$l#L       '            ����   	            ������������      ����   ����               !   #   %��������������������������������������������������������L       loss_changes[$d#L       '=���>>>��=�7?    =ʇ>�и>:�B>t�B=���            >F��>N�d    >`�    =�y/>���>�5>z�n>���>k��>�i�                                                        L       parents[$l#L       '���                                                     	   	                                                            L       right_children[$l#L       '            ����   
            ������������      ����   ����                "   $   &��������������������������������������������������������L       split_conditions[$d#L       '?�}�?:h�?�����ϻ���@n���o�?GĽC�����=ӖI��L=`��@	�F?Cн���>�`=�ۏ>^��zd�@@�=���?~�ܾ��@�I=%ڽg��;�M(�> �����=��������z=&� <�b�{=X���08L       split_indices[$l#L       '                                                                                                                                         L       
split_type[$U#L       '                                       L       sum_hessian[$d#L       'C4�C0�A C�Cv�?��@�D�@l��B�zA�@[@e@/p+@�?˙kB�k�AM��@@�A�A?�&�@�0B�x@�6]AT�@D��AYGBA�@?�a+?��4B��A;�?��P@�}�@�
7@g?\?�P�?���@���A��@�;?�]�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       39L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       G��佚";��M�WDd�L*�=.7���ץ��k���+����=���<}�~>�B�'�5;rڷ��߮���>��N�=4��V��>qĽ8�=	�� ��?u�<򃬾�X�=�]G�ז�=�⽣�g>V�<��Ⱦ�� ���s>�Ȁ�*ʴ>%�=�$ҽ��>�s���ν� _���>,�]�&)���A<a7>�f%���=�t��l˸���=�ٞ�=.��>��Ҿ�O�<��k�`-l>yս}�>��;�4�=�/>Ӳ!<�>��=&NY��M�=���L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       G                                    L       idI �L       left_children[$l#L       G               	                              ����������������      !   #   %   '��������   )   +   -   /   1   3��������   5����������������   7   9��������   ;����   =����   ?   A   C   E��������������������������������������������������������������������������������L       loss_changes[$d#L       G> w�>2l�=��=��>3@>�j>��S<�p>�o>+=�>R�?�>���>��>T�O                >dF>'z=�A�=ݶ�>�wj        =Y�/>� �>�C>�O�?J�=�:        <
E�                >���?!�        >Y!i    =��#    >���>��9>H�(>��=                                                                                L       parents[$l#L       G���                                                           	   	   
   
                                                                                             "   "   '   '   (   (   +   +   -   -   /   /   0   0   1   1   2   2L       right_children[$l#L       G               
                              ����������������       "   $   &   (��������   *   ,   .   0   2   4��������   6����������������   8   :��������   <����   >����   @   B   D   F��������������������������������������������������������������������������������L       split_conditions[$d#L       G��n�?솿R�s?cg���~~�T���L�����j?s���*�?��J�T�Z>��P>�Ӭ?���Ц��*�=?��xX�Nf���=�C@6F�)`;�F>(�_?��
�O���L�P?��x�HP=�j�;�R�� g��EW=�#ͽL�?=*���V��'V�=+���^�?�@^�Q�I���Ge?�|F��Qܾ�T�?��<ٿ��ս��}��S<Q�u=�R����;�"����=>+ͼ�I=��z�<��<�֟=��;+��>��<G�8� �-=��L       split_indices[$l#L       G                                                                                                                                                                                                                                                                   L       
split_type[$U#L       G                                                                       L       sum_hessian[$d#L       GC��A�� C��@�|Ad�By}pC��Y@\c@��A�@���Bf[c@�jA=mC���@o9?��?��@?�g�@�\�@�ޚ@+�@3B�Bb0o?�^~@��@.z6@��Q@~?gCe�lA��@5(�?�!F?��,@"E?�?�p�?ޫ�?���B'ǨAi�?�?��X@��@[=@:є?�ۧB9vIC7h�@�F�A�Z?�N?��?�
d?��B9B@h�]@*�/A>��@3��?�{l?�C�?�__A���Afc�?��C6$�@��c?�T�AR��A*~L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       71L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       =���;��
��ں=4u�~�;�Ѿt-|<���>�C6�M����$A4><I���-1=�@�=��a �;�x�qTǼ�cʾҷ�>��g�D��������"<��4>���=%g�f7>��@=R��bF>q���W"��>�v����@>�j=k���X���>� ?�w>J>���}�4�'��=
�@>�TA=��I��(�}���ܾ;>�ܒ�X|�:��a�n>Ѣ5>� �͸L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       =                               L       idI �L       left_children[$l#L       =               	         ��������            ����               !����   #   %   '����   )   +����   -   /   1����   3   5   7����   9��������   ;������������������������������������������������������������������������������������L       loss_changes[$d#L       ==��$>Ia?Hz?��?-�?!�>E{�>�.�        >�f?�P?*�l>���    ?W~�>�q�>��=��?m[    >��X>�>,�y    >ý�=Y�p    >��l>g ?=dt     =h��>�L�>�@#    >�t        >��                                                                                    L       parents[$l#L       =���                                                     
   
                                                                                                           !   !   "   "   $   $   '   'L       right_children[$l#L       =               
         ��������            ����                "����   $   &   (����   *   ,����   .   0   2����   4   6   8����   :��������   <������������������������������������������������������������������������������������L       split_conditions[$d#L       =>��о�d:�q%}��on��ƾ��j@-޾�%T>[��3*C?�N��߂�>��Ծ��<�M���i����?�˿.��>�/F���L�	в?�m�?��\�������iž55$��#P=S2?�s}<(b�@8�z�K��?A���5Tb�&*��Y�=52�������j��FE=+4>'t)=+�=����_S�Io<&E�>e�<����h��`��r$=��}�����`S���v=��s=���:��L       split_indices[$l#L       =                                                                                                                                                                                                                                 L       
split_type[$U#L       =                                                             L       sum_hessian[$d#L       =C�a�C���B�2*C�[C*"�B���A$JC
��@,b�?�]sC)�B��Ady�Au?�]C��@UBC$i[@��mBw�T@(��A4�%@>a@�]�@��.C�A@da�?�>i@��C!�:@HL?�9�@g��@��zB\΅?�2�A$��?�BO?��s@QP�?�ՖB��A�@n�?��~?�y?�2AB�$|B���?���?���@?�љ?��#@��1AFX%B+8|?�p�A��?��?���L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       61L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       ;P��x��=#��Z[��_�>V�F<���o��>��ƽ X>�7�>���;ab�^�r�R������<����c
>���=����/�Y�=������1{����<_�>^��m�)L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L                      L       idI �L       left_children[$l#L                   ����   	      ����������������         ����      ������������      ������������������������L       loss_changes[$d#L       =�t�>h� >+c>e�7    =�>>9"�>J��                >_Tt>��>�s    >7h>	�            >��>*�                        L       parents[$l#L       ���                                                                                      L       right_children[$l#L                   ����   
      ����������������         ����      ������������      ������������������������L       split_conditions[$d#L       >:	=��I��=ń�������>{a�<�f�=����@j=��R=�]�>��a:�zH������`����r>w�=�(<�Ǯ��9u>��?�$ƺ�U��T����;6�="q����L       split_indices[$l#L                                                                                                                      L       
split_type[$U#L                                    L       sum_hessian[$d#L       C��B���Bg��B���?���@zH�BXRB�p=?��?�[?@0(?�Y#BQ/�B�=X@�.L?��&BJ��B��@N�?�1@DA���A�7�B��@~��@D�<A���An��Auz�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       29L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       5�0Iݻ���=�� �K���ȓ>Oϋ=,=��O湔,>0�޻�����Q >�m�>���\������Ĭ�>�����"�_��`�>�m�=_9�>�/Խ�z|�e[�>L�ɽ��_>����Y>@�����>;a�> �&��m=�`>�P��9#{=S�����=C����/\>�<�? �#=�ҽ�:��������>@���e�b`'��f���<JL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       5                           L       idI �L       left_children[$l#L       5               	         ����      ����         ��������            !��������   #   %   '   )����   +��������   -����   /   1����������������   3����������������������������������������������������L       loss_changes[$d#L       5>��>S b=��L=}�>��=Ԁ�>�@<��    >�v�>i*�    =(Y>k�[>�tq        >��~>��>���>z3�        =a�=dZ|>�f=���    =��         =qSp    >ץ~>��                =��X                                                    L       parents[$l#L       5���                                                     	   	   
   
                                                                                 !   !   "   "   '   'L       right_children[$l#L       5               
         ����      ����         ��������             "��������   $   &   (   *����   ,��������   .����   0   2����������������   4����������������������������������������������������L       split_conditions[$d#L       5?ܭ��j��@SM?M$�f�\_?�7�m�渱�h>�*�c'�cͿX�<G.?�����Fʼ�S;��?AȾPI��]r�=��]<�2f>��J?n�X@Q8�Ѯ�>u���k=gc��:�=`�i=R$ֿ[�D<��=ߔ`�^*�<}�ʾ�H�<j�"��8=�{�>��=x����+p��!^=f��������K���Z���L       split_indices[$l#L       5                                                                                                                                                                                                   L       
split_type[$U#L       5                                                     L       sum_hessian[$d#L       5C���C�v�A�r�@��C�B=@zn�AHIc@L=�?���@�H�C�]?��@-�(@��@��H?��$?��U@��q@Zw@�(�C�\x?���?���@B��@�P@��B@0$?���@�Q?�D�?�pX@9�S?�vEAO��C��Z?�@[?��?�U�?�&�@Ny�?�Y�?�W?��@&��?�??�d`?��F?��^A<�e@�?C�A?�vJ?�}5L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       53L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       +�'9;0�W��U�:4u�>8�u�E����!B>w����=#��>�s�<�FN��V�>D
\��o^�;d*>z�!�-�����¾����Ct¾��p:Pf�>�T���C>�\��3�=�~?��l�>|��O�ɽ��=����W�<��>���=(���V��u�¾�ux=��E>�[��@�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       +                      L       idI �L       left_children[$l#L       +               	            ������������   ����               ������������   ����   !����������������   #   %   '   )����������������������������������������L       loss_changes[$d#L       +=�aq>�-=���>�C=>t=�d�>��>u=��            =/v�    >�K=�ʹ>��>R�6>��\            =�u�    =9�h                =��>h�K>��`>��                                        L       parents[$l#L       +���                                                                                                                                  L       right_children[$l#L       +               
            ������������   ����               ������������    ����   "����������������   $   &   (   *����������������������������������������L       split_conditions[$d#L       +?ܭ�?�C�@SM��[O?��޿\_@�b�?��y>�<D^a=��<����V=k?���=�o3<>�L@�҉��i�U��e�j���0 ?�7=W2�m��> ���=���=�ʿf��<G.?�U�"�� �;�
�=���<I����4ݹ�Y۽���=T�=�n�f{�L       split_indices[$l#L       +                                                                                                                                                           L       
split_type[$U#L       +                                           L       sum_hessian[$d#L       +CƮAC���A�JoC��`@QR@q<BAFE�@�ZC�)�?��?�'�?���@$��?��RA1σ@{ߡ@j�x@L��C���?��?���@
]�A8?�z�@�F@9e?�6&?��)@�Q@N�nC��y@�/#@�@�?���?���@
��?�.?�l�C� ?��O@�@87�?���L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       43L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       O;+�>��&<�79�^6Z=x�t~=���Ŵ=,>.ĝ����yR,���>E�<�L�_Q�1?C>u⣾I�>��=V������=�`$�i"�>U�ݾ���U��>��D��n�%ؖ=j�>=�o�K�����	<к->�]����l���.=�΄��C�>3�U�']�>%�[>�Ǭ�U�����#>�o>�J�=��7�s^;=>mm ����j�>S�¾��˶�[Q��Vҽ(�;>����ب>�U�=Z}m>XY��)��Z��=��4>��ʼf9`��F0����= �����=���H�<>�Ť��L��b�X<U�TL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       O                                        L       idI �L       left_children[$l#L       O               	                                    !   #   %����   '   )   +   -������������   /����   1   3   5   7   9   ;   =��������   ?��������   A����   C����   E������������   G   I   K   M��������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       O=�e�=�<>�>D�>0�C>\G�>>�>,/>�h'==Ќ>��>9��=?%`>��V>'��>���>��F>Y�4>�2?    =���>:$>���=��            <t�@    >�*?0J>r�>�=;>��D=���        =���        =�d�    >z"    >�            >�X>�>.d>�R                                                                                                        L       parents[$l#L       O���                                                           	   	   
   
                                                                                                           !   !   "   "   #   #   &   &   )   )   +   +   -   -   1   1   2   2   3   3   4   4L       right_children[$l#L       O               
                                     "   $   &����   (   *   ,   .������������   0����   2   4   6   8   :   <   >��������   @��������   B����   D����   F������������   H   J   L   N��������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       O��8?���:R�>�O���[P�H�!�(f���m��C!��׮�@	~��XCe�pp�m���1㠿$Rڼ��I���o=��?�1�L?��g��R:�Q��=�R�ޛ㼀V)�mw�$&��U�ǮO�I7>El���nD����(�R��>���?I�T�(�=W� >��h=F�n@����b��g<@=,��=��5<�^��q�\�(��?��a0���=}��ʭ[������4��J�{=�(@�8��=�3�<�=��ϼ�˥��]H<Ћ>����"m�÷����<=�ս��<�/8�p�|=� _��[����h;�f L       split_indices[$l#L       O                                                                                                                                                                                                                                                                                           L       
split_type[$U#L       O                                                                               L       sum_hessian[$d#L       OCj�B[��B��lB�|A���A�<�B��=A���A@��@�iMA@�A`3�@!�@��?B�yAO�ZAN�@�j@�a�@�u@1%Ab@^�A<�A@�E?�#�?�>@Cz�?��nA��;BK"UA W@�v@�D�@��r@zQ?�a@?�@s�/?�ӗ?�N�@�a?�[@G�?�ƙA"|�?Ѻ6?��?���@�7�A��UA?�(B2@dr7@�Œ@%�@��@�݆?���?�@PR[@2�u?�m-?��@�p@�y?��(?��?��OA\f?��?���@�]A��K?�P�A/�?�S�?���BZ�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       79L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       �S��On:� �I��<���!;�Ȿ|���#d��:K=���>1<�;�S=y�^_Q>t��FJ-�g��;n䅾�0н5�/>�A�<Q��>���;���gI=.��N��<���L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L                      L       idI �L       left_children[$l#L                   ����   	   ��������   ����      ����      ��������   ����   ������������   ����������������L       loss_changes[$d#L       =��:=J�x=ЦI<�[�    =č�>��        >��    =��=�>�    =�:�=�L�        >]�    <�:�            =�                L       parents[$l#L       ���                                         	   	                                          L       right_children[$l#L                   ����   
   ��������   ����      ����      ��������   ����   ������������   ����������������L       split_conditions[$d#L       �M��?��;�8\?sB�;73�?��;��������DG��D�<��?fǾ��3<�ro���V>AA�m򝽊虾��n����?��?=߂;{p�=���>;Ƚq,<;k�xq;ؼL       split_indices[$l#L                                                                                                              L       
split_type[$U#L                                    L       sum_hessian[$d#L       C��w@�C��#@OW�?���A
	oC�1�@�,?��@�	0?�&�@�l�C� $?��(@�J�@HN7?�?�r�C�u�@:#�@qf?���?���?�p�C��A?��?��8C=��C
H�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       29L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       ����;�P���z9s�
>�[��h=�_�;�l�&�>��S#s�"�>���:Y�>j�^>:-���l<IY>f����྽o�`;*�C��&t=�#���r&���>:�P>`�\�ځ�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L                      L       idI �L       left_children[$l#L                   ����   	               ��������   ������������������������      ����   ��������������������L       loss_changes[$d#L       =��I>C�)=���>J    >���>J>d>�d>��/<�H>=a�        >.�                        >%K�>U�q    >�                    L       parents[$l#L       ���                                                     	   	   
   
                        L       right_children[$l#L                   ����   
               ��������   ������������������������      ����   ��������������������L       split_conditions[$d#L       ?_�?T?�*F?;B=��>3�?��?7�����ƾo��?� �C^�=�%�?-M�=���=_j���;q�!=�p���~?Q�?����.%�o�콡Uȹ�=`Z�=����L       split_indices[$l#L                                                                                                                    L       
split_type[$U#L                                    L       sum_hessian[$d#L       C��C�U�AE<tC�j-?�<AN@+�oC�_@���@	�@�a?�2�?�@WC��.?��;?���@.�W?���?�UT@54�@�s�C���?�Yd@T|�?���C��@�ј?��j?��L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       29L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       /:�4�,��=���<�:J��n#�i�^>p�W<0�>B�����E=O">�}��&ݼKh=�5">�nf�������&=���>f�.��nN��P��j�;���>����Ҷ>�>(�V�F�>���<��=)��4���3<�<=�l�^��>���=��{�F�h�$�k=[��>��[�*�/>�ھ��ǆ�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       /                        L       idI �L       left_children[$l#L       /               	����               ��������      ��������               !����   #   %   '����   )������������   +   -��������������������������������������������������������L       loss_changes[$d#L       /=�gi=��.=�z>QR>-     =�̎=�->�>7�>P�        =��c>U�,        >r>=�L>���=�ZG    > ��<��=�h,    =,��            >��=���                                                        L       parents[$l#L       /���                                                     	   	   
   
                                                                                L       right_children[$l#L       /               
����               ��������      ��������                "����   $   &   (����   *������������   ,   .��������������������������������������������������������L       split_conditions[$d#L       /@*It�d���L.?K�?�9��Q����d����~?��?�t=�60���=>�ȿ?��=��{��n�@@W�@3	6���?dk�W�0����H�^�A�E>b8R=/Q2>B=�.U=��m;�?��?�` �˙;�H<�������=�#�<����n�}�E�<��\=���M9=����g���n]L       split_indices[$l#L       /                                                                                                                                                                           L       
split_type[$U#L       /                                               L       sum_hessian[$d#L       /C�C��@�B�B��eB���?��@BB��)@���B7�A���?��'?�I]Bn�A)U@<�?��B1@� �@n�(A�:Bj�`?��@��@A�Bb�?��*@�!�?�}6?��?�cA��@"�AF�rB9�@�F?��h?��?��0A�B�A��I@2�?���A�A	��?�P?���L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       47L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       ;������6�;��X�Ԗm>/89A��=�~\�A!����]�AZ;K�=&�>����H_���jo>A=*���������W>-H���Vy=�$��辐4k=����n��0e=^�>��A<��:�T&-�
T=�^�>������u�N^�:�ꢼ�0>P�	>j�s��콂��>x:��m>ᾚݐ�T�,��Q>��澘�>����R>=��;�mݾ �d>	�o�/(}�N$>�g�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       ;                              L       idI �L       left_children[$l#L       ;            ����   	                  ����               ����   !   #   %   '����   )����������������   +   -��������   /   1   3   5   7   9��������������������������������������������������������������������������������L       loss_changes[$d#L       ;=��>$;=��Q>%B    >1��=��{=�Ѵ>]��=�@�>v�>�
    >@!a=�CD<�cP=�wJ=���    >���>G��>/r?ݠ    =�v�                =o�=+2�        >wP>F��>�1�>A?>H�>1U�                                                                                L       parents[$l#L       ;���                                                     	   	   
   
                                                                                 !   !   "   "   #   #   $   $   %   %   &   &L       right_children[$l#L       ;            ����   
                  ����                ����   "   $   &   (����   *����������������   ,   .��������   0   2   4   6   8   :��������������������������������������������������������������������������������L       split_conditions[$d#L       ;��n@\~?ܭ��|��=RCT�j���3�L�*�?�N�m�l�fؾ�H�=�]��N�4<��]>#�Y�����n޲�Ѷ>�*�c'�@�\?��ܽ���N߽ډ���z<*�:=��N�����R�%�2=8�;ҟ�?4�:�PI�?βH@�T�z=��E�����&�=�﫼ٶ=&꨽�֭���aB=���R�=,cͽ�|c=cnU:�P��A$=%b�R0���,=�|�L       split_indices[$l#L       ;                                                                                                                                                                                                                         L       
split_type[$U#L       ;                                                           L       sum_hessian[$d#L       ;C�Y�A�C��'A�!�?�X�C���A{l0AB�A
@q��C��Aa�?��@��@���@3�@�"@y�?�u@��C�]�A;��@�?�;�@M,@f�[?�v?�8�?�G_@+� @8�?�IQ?��i@���@�@si`C�v�@�T�@��*?���?���?�,�?�+^?���?�Y?��?מ?��Q@���?�%�?�~W@1�?�b�C�Q�@�U�@F��@S�	?���@Y��L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       59L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       )��(;	 �����;������Z=�����;iP >)���2��И<0T��@SN=� K9}��=�>��Ľ��3>6{T��>B��N�<��>�|}���p; L<��߾PL�VJ�?���܇>,=�z�
�]>��H=��i=��C�<�y�	Jq>0R=����I�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       )                     L       idI �L       left_children[$l#L       )               	����            ��������         ��������         ����      !����   #   %   '��������������������������������������������������������L       loss_changes[$d#L       )=�_I=�3}>`=��>�    =x�(=ǫ=�`>5�        >!>)��>@�        >0�?�=���    >;��9͐     =�_�>H�{>1{�                                                        L       parents[$l#L       )���                                                     	   	                                                                  L       right_children[$l#L       )               
����            ��������         ��������         ����       "����   $   &   (��������������������������������������������������������L       split_conditions[$d#L       )?� ?ܭ��h�?�C��3�L=�߿���i�U?��޾�H���-�;S����@�r���f��<>�v=���@�\?��ܾ��ƽ��ǿ�[O�W�ƽ����`ن@�T�z���N>'%�$;�=-�=:��&j�=ğ�<�j�<�y�b���$��=SJc< U���X�L       split_indices[$l#L       )                                                                                                                                                     L       
split_type[$U#L       )                                         L       sum_hessian[$d#L       )C�aC�giAC��TAr�?���@� DC�4�@M��A^w�?�V�?�K�@�mVAW�C�w�?�=m?�xFA;^=@f@2�r@<W:A0Ű@]I?�(PC���@�@��_?���?��^?���?�:@�}�@r?�k]?�O4A�VyC��&@F}�@S�H?�̽@Yv_L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       41L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       Q;(B�s��=0�L��ڕt=mY#��M����=�l�Z��=n�b>���v;< �����X��$�<Rq�o[O>i[�=xBz��_�>�������-��>Q���X>N'��[�=�O>O�N���>W�T�������s�1^;;�X�>�J���=x�3D��`ǌ=�j=V�=�_�>�O~���=���Gc�>�]=�U���=��>�q˾���$�>�������|��=�[%>��xq�<���>��=T��.�R>Z�u�wgD>�����.>`��^g>4P=��*����=�Ȩ��`�>F����>�nV=;�m=���>(L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       Q                                         L       idI �L       left_children[$l#L       Q               	                           ����         !   #����   %����   '   )   +   -   /   1   3   5   7   9   ;������������   =����������������   ?����   A   C   E   G��������   I   K   M   O����������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       Q=�3=�2�=��"=��M>M�m>��>
>��?�>>(�t>nod>fcR>m��>$�k    >�J�>�m�=��=��t    =vY    =�Uh=��K>�q�>Mb�<���>��>�u>A�~>玦=�X>��|            >"�p                >	��    >GRH>�2J=��q> ��        >�̈=:d>$�>�                                                                                                                L       parents[$l#L       Q���                                                           	   	   
   
                                                                                                                       $   $   )   )   +   +   ,   ,   -   -   .   .   1   1   2   2   3   3   4   4L       right_children[$l#L       Q               
                           ����          "   $����   &����   (   *   ,   .   0   2   4   6   8   :   <������������   >����������������   @����   B   D   F   H��������   J   L   N   P����������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       Q�K�l>z�?��<lgA@	���M�V@c�6q�:�¾�@�@=ؿ?��@�9?8L���7�!�0��^�Db翓&<���@�=���@O��H+U?6\�=+�?b�?�?�Mp�E�t���H���`�gŹ��)W�T�{;5c�F� ����W����!<�e��X)j�����4?��?����RV=�<�<=y��N�?�f�>�Q�?���Ȓ�=�P"���J����<�m`=�&C��1;�G�=��f<~}�Q�=�)z��q)=��3���=�sr�8
�=X`<�g ���J=����y=nvm����=�<aN�<�P����0L       split_indices[$l#L       Q                                                                                                                                                                                                                                                                                                    L       
split_type[$U#L       Q                                                                                 L       sum_hessian[$d#L       QCb�B��BW�&B��MA�nBC8A��B�_�A�@�e�@�A��'A��IAp��?�P�A�BF��@%}�@�k?�l@�a$?��Q@ ��A��AQ$�A`�@�@���@�|v@&ޚA�C@@���B/��?�m?���?ݡ`@��@N��?�v�?�5^?��@�]%?�(�A$\@3"<@޺�@�b�?��?��@�!@m�C@��:@-�v?��N?�8�@пAv&�@@j�@1b�@��B�@>(b@�-@���@��?�A�AS�?��w?�S @���?��?� 5@���?�ҷ@<��?��?��@��@��?�6?�6�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       81L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       5�}�ʼ<��<瑤�e�&�78��y�=P�|��p=���>��ҼDxh�[�=�S���J=��¾<B��o�=�������><��=��Q�B�->���=G��>w�ھ�`�>kV�]t5��:x�{&=��?���n>x鑽������>��<�1>�L<�\�>F?۾�w�>��H�R縻�Ā>JV��+��2L:]"(=K徳!P��>�WL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       5                           L       idI �L       left_children[$l#L       5               	      ������������                     ����      ����   !   #   %   '��������   )   +��������   -������������   /������������   1   3������������������������������������������������L       loss_changes[$d#L       5=ڒ�>@kJ>��t>=��>��w>u��>~            >I��>nZ>=��>mE�>�T?*��>b�?    =�'�>�i    >	�">���>'R�>��         ?H>���        =:
K            >D��            >�K>��                                                L       parents[$l#L       5���                                               
   
                                                                                             #   #   '   '   (   (L       right_children[$l#L       5               
      ������������                     ����       ����   "   $   &   (��������   *   ,��������   .������������   0������������   2   4������������������������������������������������L       split_conditions[$d#L       5>��пh"�>mf#?F�^�f�u��G��؆l<��[=��c�^sпK��>ī�ij��=Vp=�6��Y^<�#S?]yL=�2=bL;>�O��Om�=sy�>�=����s�?�?�T����F*�6�.?�g���QQ=�X���?m/=6�<�>ka>��F�0S<��)_=��$�}��==�μ�A� ��9��<:[���ǽ �=���L       split_indices[$l#L       5                                                                                                                                                                                                  L       
split_type[$U#L       5                                                     L       sum_hessian[$d#L       5C�IC}p�B��>@E�Cz\yA^�5B���@�?��@  �Cx[�@�2�@�U�A�uB�<I@��&Cr�6?��@��}@��?��2@K3�@��@�b�B|L5?�y�@o��A��Ci�@v��?��Y@�n2?�ש?�Ն?��a@�8�?�O�?�/�@2-�BQp�A+n�?�\�@�k�@�/Cc�k@!?ӊ�@Y�?���BI�@�@,ӒA 9�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       53L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       E��Ֆ;��E�)Ɉ<���.����=T�;��>����D�i=��T��n���=��н��?;��>�ɾ�H�=�wu>A���B$�<�3�����>b�
�I;�=1�þ�r���B�=�C�:sL>�5w=�R��N�0m>̜���<>�-&����;ug>������P�Z�>��>����l�;�2��۹�>�V�<�0��b�<�g >��=�^Ὕ>��~p=��P��N�>҈=�!H���1��x�?��=�\����>V.����;���	>���L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       E                                   L       idI �L       left_children[$l#L       E               	         ����         ����               ����   !����   #   %   '   )   +����   -   /   1   3����   5��������   7   9   ;����   =   ?   A��������   C������������������������������������������������������������������������������������������������L       loss_changes[$d#L       E=��8>�f>��>ae�>i��>���>��>)     >�<>S	Y>�:�    >�#>�dG>�C?ȸ>F�*    >�     ?�K=�;�>�p�>�a">!|�    >���>��h=�v=�P�    =p        >���<��=��x    >�a=��(=�9|        >��y                                                                                                L       parents[$l#L       E���                                                     	   	   
   
                                                                                                           #   #   $   $   %   %   '   '   (   (   )   )   ,   ,L       right_children[$l#L       E               
         ����         ����                ����   "����   $   &   (   *   ,����   .   0   2   4����   6��������   8   :   <����   >   @   B��������   D������������������������������������������������������������������������������������������������L       split_conditions[$d#L       E?|�G@�"��j@
pw@@�h���!��M�?z��=�k�>AA���1i� Y5?���H�J?���>l����'<����)��h���O�	>������@5���I�(���?�� ?ڣ���?���<�b�Li�S�%=��˿a��?;�>�h :�>?�GV@ ��@S�=�f�=�n��:�<����=��@;.���2;��>��<�>������d�<�����+�=��F<�[$������Q>$�<�o,�,S=)����Q�:�
��$h�=���L       split_indices[$l#L       E                                                                                                                                                                                                                                                           L       
split_type[$U#L       E                                                                     L       sum_hessian[$d#L       EC���C��8B0�+C���AAT�A�AԧRC�f?�+@�r}@�7[Aw��@	��As0�A6�C�3Z@���@�9�?��@W�?��A'/@��A�@���A	�@4W�C�	�A��'@��@^��?��;@�J�?��^@��@�F@*00@}??���@��~@f}I@uy?�p�?���@��C�A���@�{�AonT?�4?�)�@P?��?��@vF@��G@VZ ?��?�x�@6i�?���@L�E@0��@"{?�ɜ@l�?��@���?��L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       69L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       =;F_��u�<�Bľ&�+�޻���=��-=9`4����>�UL����<�)�e��>b��<����M:"<���<�:ͽ�(�>�$p=P�z�5E�=�����(Q=��>�ռ�$���~�=� ,<��C7�=fl�>ĺ����=�ի>�&�߽����<�F>h����f�>q'V=�ӽ�=���=���=�)>`�3�l�h=Զ�������Jo�Ṋ=��Y>7X���=�k�G>=�{�����5YCL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       =                               L       idI �L       left_children[$l#L       =               	      ������������      ����                     ����   !   #   %   '   )   +   -   /   1   3��������   5   7   9   ;������������������������������������������������������������������������������������������������L       loss_changes[$d#L       ==�%M=�D=޿>a�>#�7>K�>cV�            =��6>�z    =M�0=���=�f>P�>�=�|Q=�V`    >�P>�=���>��X=:��>z�>��g>�>�<ѿ==g�@        >!4>��>��<��h                                                                                                L       parents[$l#L       =���                                               
   
                                                                                                               !   !   "   "   #   #   $   $L       right_children[$l#L       =               
      ������������      ����                      ����   "   $   &   (   *   ,   .   0   2   4��������   6   8   :   <������������������������������������������������������������������������������������������������L       split_conditions[$d#L       =��8�w���1������it���à�QB<^sr��ra=�3(?����(z���(<�����J>ѯ���[P��V�=���%[�<z��?�{x>�o>Fz:�C!��׮�>	��(�4?�r$?A4�?��<�AQ=�'?q�?
����_4>����+��;��=����
h=��4<;1��}7=a^</�սc}e=<ٶ�'
����<�A����պ򿹽x(�=i=\��㼍c�=c�������Y�QL       split_indices[$l#L       =                                                                                                                                                                                                                          L       
split_type[$U#L       =                                                             L       sum_hessian[$d#L       =C�BRœB�Ch@��OB?�)Bp��A��?���@6��?�'8B;H�Be5�@8~�@�9^A��A���A��_BM�b@���@���?���A;�#A`fgA�7�A ��@�A5�A��A���@�:@y��?�r�@�S@�l@�0�A4J]@0p&Ai��@���@�j@� �@
{�@%�sA�@C�%A�;@@��A���@��M?��?��h@&�y?�n�@�h?�4@S�?ړ�@.��A��?�%�?���L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       61L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       -��m���:�:�����=�.>F�Ǻw7�y�;Y>�>��ռ	Xr���;_�%<9H���Jk�"�=�J��s�)�~\<HOh���Z>!K�������C��cz���z=�g`;��.>��վDȋ<���$�<��`;d����M�>{>߽��<��Ⱦ:�;$[�>�������6��&ad=��9L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       -                       L       idI �L       left_children[$l#L       -            ����   	         ��������      ������������               ������������      !   #   %   '   )   +��������������������������������������������������������L       loss_changes[$d#L       -=�d�=���>��>
;    =ҥ =ߚw>�V=���        >E�=��            = Ϛ=O�@>#!�?'Z?T�            <��F>y�=�ti?s>U\l>��F>�;                                                        L       parents[$l#L       -���                                                                                                                                      L       right_children[$l#L       -            ����   
         ��������      ������������               ������������       "   $   &   (   *   ,��������������������������������������������������������L       split_conditions[$d#L       -����?�o�����>U��<�GѾR~���n��z>�ŵ=����$Љ�@Vۼ�l";^W���&�B�y?x<�?RP<��a���>��w=A���Eӽ�Ʉ�C��Ï?��J>��>��/>~�h�D�_;�+�:�.���*J=��S�/;�y��`O:E:�>���,�*�ܽG�<���L       split_indices[$l#L       -                                                                                                                                                               L       
split_type[$U#L       -                                             L       sum_hessian[$d#L       -C�ǬA�yC��@�|�?�'�@HӐC���@��k@s�?�p?���A���C�!J?�>@0��?�!�@/VA@�#�AICv�B}
?��m?�?��@?@@�%�@�ޅCs �@��A`�BDυ?�R�?�+�@�l@"�@�<@��Ce֜AR�h?��.@3�AKB�?��A*1BC@L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       45L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       /9n�ܽ��?;/��>9��	��=ǚ��(��H�A=ԋ(>$hk���޾Idi8�P���羬�����\>���=���Zs�<�N����>t��ֳO�U��>b�=�ݪ�,c�>�~�<�»��I>$���ڋ�5�Ž�:;�������26>�ݎ�7SP<xH���	D>�9.=��������>��=�W�sL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       /                        L       idI �L       left_children[$l#L       /         ����      	      ����               ����            ������������   !   #����   %   '   )��������������������   +   -������������������������������������������������L       loss_changes[$d#L       /=���>?>?m    >,��>h>:T=�|    >�Ų>$=��|>��>���    >+�+=��8<�ß=��            =��g=�ь    >�5=s �=�I�                    >��>�9                                                L       parents[$l#L       /���                                               	   	   
   
                                                                           !   !   "   "L       right_children[$l#L       /         ����      
      ����               ����             ������������   "   $����   &   (   *��������������������   ,   .������������������������������������������������L       split_conditions[$d#L       /��#V�oͿ`�=_$ܾot�=�Kj�Vix�C<�d�s�C�;�H���Tva�!����|��R��מݿ]{�Ҁ<bf��K�=�n��g�D�g��=��ʿ~��!�;�l�<註d,=D�ͽğۻZ@�g�P��"�����<A=�=�[��;��k����=��8<��ڻ��7�,�=�氷�\�L       split_indices[$l#L       /                                                                                                                                                                              L       
split_type[$U#L       /                                               L       sum_hessian[$d#L       /C�^	A'#*C�$�?�KBA��A��rC��@�p?��OA\@�ɞ@p��C���@��@?�ܿ@�c@��@��@%�H?��k@&��?��wC�'K@�,B?�G�@�b�@']z@�_�?��J?�a�?��J?�w�?�p�Av��C�q�@Gr�?��n@"|�?��h?��?��@�/�?��PA_��?��7?�NC��gL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       47L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       I;5F����=H�<��p�M��=�F���:���=�=��
���g>M�P�J����L=�<!<.3�(%L>�Ť=�޾-�=��>�W���=]�Z>�%����=�p�j�>ִ>�`�����9>R�Ⱦ�He=���;蹼>\Y����H�O|>�y�=�AE>\$ľ�'>�V�<��#>ɽJ�%��(�=��>ǫ�<���?�p�E$�<.*�.�>���<�RU�ܦ����^�%�Y=�K>����#�̾IN�>�|�p��<���=I�ϽYd�<Lq_>F���,���L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       I                                     L       idI �L       left_children[$l#L       I               	                                    !����   #   %��������   '   )   +����   -   /����   1   3   5   7   9����   ;   =   ?   A����   C����������������   E����   G����������������������������������������������������������������������������������������������������L       loss_changes[$d#L       I=�u>n�=�r�>߰>I6�>���>Q�>&�+=�� =�d>C�p>~>g�>G�>��^>�r>@Q�    >1 =m/X        >&�>R�b>C�d    =Vli>/c�    >�h<Ճ�=�a�={G�<��    >fS�>Ձ>�=��     =���                <ߙT    =�j�                                                                                                    L       parents[$l#L       I���                                                           	   	   
   
                                                                                                           !   !   #   #   $   $   %   %   &   &   (   (   -   -   /   /L       right_children[$l#L       I               
                                     "����   $   &��������   (   *   ,����   .   0����   2   4   6   8   :����   <   >   @   B����   D����������������   F����   H����������������������������������������������������������������������������������������������������L       split_conditions[$d#L       I?GĿd�?��:�zH=��E>�,?8L�����v@UT>�?�Ɓ>�Ol@`]?�T�?[/D�� g=��žy����<��n=�����e�Z|(?������?��S�8z�=4ؾ7�V@�}?b��?ƃ�U_�<�f>:	?�*u�ފ?������>xn=��6�> �o;�:������s`?<4K<��=�;��:�fT�l��;P�f�PԠ=���;�/��c�щ��F��<�i'=�&�DP��q��=*L����&;֜�<r���o�;uT�=n�%�7'Ͻ���L       split_indices[$l#L       I                                                                                                                                                                                                                                                                        L       
split_type[$U#L       I                                                                         L       sum_hessian[$d#L       ICL�B�mSAܱ�B�F�B0L�A��A5&�BU��A�$AATZ5A�l�A� @�h @�e�@���BB@�D?�~A��YAD.??�_�?���A�|�@� @��@:�@�J�@�0�?��I@Q�@
�B7.�@.Ci@P$�?��3AH9,@c~@%��A�N@�=A��@�h?��1@G��?�4s@G�?�֖@\�{?��?ټ?�IN?�� ?�� B*��@H�f?���?��0?���?�iN@��A-^@�?��?�?�9{Ah?��NAb�AWx�?�|�?��t?�í@��L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       73L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       5��\��	;ݾ?�5�T1:?`>[����o���=�3��Ϥ�=�0���`������r̽Q�n>lU���<O=M��<b׽>��.�g:��>=�/)���=,�+>��󽘮�>X=����an�<�Np?w'��*=��>w����p=,,��wc���=�=,�>P�K��ӎ>g#�=8ex�������|��t�>q Ͻ��ԾE��;%��L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       5                           L       idI �L       left_children[$l#L       5               	   ����   ����            ��������      ����            !   #����   %��������   '   )   +   -��������   /   1����   3����������������������������������������������������������������L       loss_changes[$d#L       5=���=���=��K=f?h=���=�i�    :��     >#E�>�Q">��>�P�        =��S=\�p    =���>]�<>'r�>ob>?��    =�;�        <�pB<#�8>�g�?!>�        >ip�>
h    >Y�                                                                L       parents[$l#L       5���                                               	   	   
   
                                                                                       !   !   "   "   $   $L       right_children[$l#L       5               
   ����   ����            ��������      ����             "   $����   &��������   (   *   ,   .��������   0   2����   4����������������������������������������������������������������L       split_conditions[$d#L       5��n�?�@7��?�8V>Ϫ��R�s=���?�a���,>�?m�$�S|��L�����:��V����8?��|��{���K?�7?���>�Ӭ�K�=������<O�=�c$?|�K=�O��Z�Q�Z�2;�^!>[ɿO��?�Z�=��<�F�H<N�뽔n��7Kk<�<O`	=z�'��dE=��#<]F�������j���=��I���e�m�:F�L       split_indices[$l#L       5                                                                                                                                                                                                   L       
split_type[$U#L       5                                                     L       sum_hessian[$d#L       5C��WA�1C��E@��(AR�C�g�?�r0@HK�?���@λ|@�c�Bl�2C��m?�>�?�Y @t*�@)L@�@���Bb�2@o�A1�Cx��?�,�@%a?��?���@V`@Y<A�eyA�R�?��?�	�@��@_0@�KCvm�?��'?�|�?���?�$?���?���A���A1��A�^'@��@�9@P��?��/@�@���Cq��L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       53L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       3:
p;98���_c<\;���+{�=���;p�U>�����V#�͐�*���u5O����=��=���>�-�=��y��0>7S^�~�]�7��>�����m���b:�m���=>KP���UQ�\x�d�>����,J�`X����Ļ(/>����0��Ox>�B�yx��G�=괍>ƣ!��o�>2�ҾN�>��M�)�=�Ⱦ�]LL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       3                          L       idI �L       left_children[$l#L       3               	   ����                        ������������         !����������������   #   %   '   )��������   +   -   /   1����������������������������������������������������������������L       loss_changes[$d#L       3=���=��>o~?$}>�=Q^    >�{<�� >�g�?�> ��=XQ�?27!>�V            <=� >��>��                ?~g=&L�>���>���        >��x>>!�>�;�>A��                                                                L       parents[$l#L       3���                                                     	   	   
   
                                                                                   !   !   "   "L       right_children[$l#L       3               
   ����                        ������������          "����������������   $   &   (   *��������   ,   .   0   2����������������������������������������������������������������L       split_conditions[$d#L       3?
�>"��>���=�&W>E����X<����)!z�^ �i��gJH?��?�����?��Q=T�>N�=%�LN?;\�=���\w=;��ֻP��Hܾ����i���[�>�ŵ�';Ľ-E�?���x>�]Z�ݑ��I� > �����	�=�jP��g⽛"�=һ=�][��=VIɽw=l=Ʈ]�K��<7�ӣ)L       split_indices[$l#L       3                                                                                                                                                                                         L       
split_type[$U#L       3                                                   L       sum_hessian[$d#L       3C���C�>x@�C��Bb��@�S?�G C��D@�Y @m��BS�W@*ښ@E<C��8A� �?�u�@�?�+@$_aA2��B&�6?��?���?�ͩ@�8C���@u�@A{�[AR?Ƃ�?�<@��@ed?B2Y@�f�C���?��?��X@$�A@+[@n @��Y@���@�*g@
��?�"%@�-?��7Bڰ?��@��L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       51L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       ?:���g�=	T=�U���O�>V��<�W�����>h����7��S>���=s��6�>z>X�|�r=H}�>�ɸ<[�;�=ו>��hA=x�2�+�O>��<�h�>�����Nh��E=ٝ���>=���G9>Tu��-r;�1l�:`=��O<�{i�ϥ�Hǡ>s9>�[�>��i���μ�+�>U]���U�=�y>�w��ü���<���=&l��sK=KG>+~�<�]>9�h��,���ɻ�aL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       ?                                L       idI �L       left_children[$l#L       ?               	                  ��������      ������������            !   #   %   '����   )������������   +   -   /����   1   3   5   7   9   ;   =����������������������������������������������������������������������������������������L       loss_changes[$d#L       ?=���=�,>
�>Wi�>
��<c�0=��#>Kfd<�+@>|�@>$>�        =Խ$>S;            =��@>ꄽ>�ܲ>H>`�x>���>�-    >���            >�Uj>j�=�\    >�>�=b>,Z�=��K=p�<=�͢>��Q                                                                                        L       parents[$l#L       ?���                                                           	   	   
   
                                                                                   "   "   #   #   $   $   %   %   &   &   '   '   (   (L       right_children[$l#L       ?               
                  ��������      ������������             "   $   &   (����   *������������   ,   .   0����   2   4   6   8   :   <   >����������������������������������������������������������������������������������������L       split_conditions[$d#L       ?>v�P��'\?� �g�`�$Ŀ��@�f�nS�� g�����m=�H�<�:�=Ox�?�A=#Rн��<p�˿��ֿF��>�X�����gPʿ���_]=�f��=׵?��^��= ��~>^�:�ݽ�V�O�c�Y�@eӿqx>ˢ��e�{?��2�p�=��&��p=�T~���^���
=��3n<+�=��~��+�;�e:�b�齮�Z<''"=M�1;Ӣ�=^�}��i�ɖ�L       split_indices[$l#L       ?                                                                                                                                                                                                                                  L       
split_type[$U#L       ?                                                               L       sum_hessian[$d#L       ?C	�B� %B>'�@�L.B�[b@<�B2X�@h��@�;A���Bs�]?��?�	;B@��$?�u?쪴?���@JA�AA��A:e�@�(�BZ�IAoY�A�U>?��`@^��@��?���@ 5jA!��A�@5��?��@��8@�إB>84@#u�AF|�Ap��A�?�«?٪�@Ƈ-@y@�g�?�w�?Ԫ�?�j�@@9E@�+?�@��B1��@J֊?�1�?��0@���@�t@ 6*AH�r@B��@ր�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       63L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       7�s��;p�<����7��<m�<z��>�D�g|��|�?���'L<�D�ڋ5�.m�>i�D��՘>�m�?JX�=��6��<�ػ���=ԘJ��pؾ��<>�1�����ɼ��>f���h�;�X5��z>~�<5^�"#>�D�>m?*@?��ӑ>��Y�;������b�2>�d�>���M���8A:���G��=���>����������=���L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       7                            L       idI �L       left_children[$l#L       7               	   ����               ����         ����������������         !   #����   %   '   )   +   -   /   1����   3   5��������������������������������������������������������������������������������L       loss_changes[$d#L       7=���>P�>��;?[?P?��Y>�b�    ?Jv�?���>��$?g�>��)    >�� >�x�?��                >��>�b�>ɻR>��j    >��?3��=��`>��8?MKH>�M�>�dS    >�J?|~g                                                                                L       parents[$l#L       7���                                                     	   	   
   
                                                                                             !   !   "   "L       right_children[$l#L       7               
   ����               ����         ����������������          "   $����   &   (   *   ,   .   0   2����   4   6��������������������������������������������������������������������������������L       split_conditions[$d#L       7>���z��@=1���`�h(e@5��=Ӆ��b?v�ľV6���>=W�� S������=?�Z8=��&>r��<ݣ۽�gi���>@X?�J��
6�-X��������N6>Z���_��L�>
P���,%?�3�?$ְ�B�m=���=1�>LM��1=��8�3X��B罈.�=�E�=�8��î��9�K�o�/<��=ַ.��	$��<=MUL       split_indices[$l#L       7                                                                                                                                                                                                       L       
split_type[$U#L       7                                                       L       sum_hessian[$d#L       7C�^NCig�Bʩ�B�M�C��B��?���B�r7A�n�@-�`C
)B��?��|B�H�A9J�Af�<@dd?��?�/;@#B���B��A�PB�%@7�@�5�@�_�A",�@���@�خB��.B�B�?���A'}�A�U{B��@��@�k@��?�=T@��@��G@�e�@A��?��~@�`�?���?�׿B��B��A�KU@��@E� @CҧAo�ML       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       55L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       ?8��R;K諽�?<�v��-� 4�=̓�<�r�a!�1~=
c=A˂�TrZ��}>V�<���>�"�	(��<"���X�ę�>.����ė�=����Z��-��=��#�hRټ �>���<ր����½�þ�o>�gɽOՅ�W?>�Z>)}�<�΃���M��K<>}Y�TD�<�#~>��/��`<���<(�ֽ�S^���>�����9W{=�@�>�l��	�"=��0���ǭ�>���D�eL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       ?                                L       idI �L       left_children[$l#L       ?               	                        ��������   ��������         !   #   %����   '   )   +   -   /   1����   3   5��������   7   9   ;   =������������������������������������������������������������������������������������������������L       loss_changes[$d#L       ?=�>�=�)U=�+t=�і>�.>-�
=���>��?n�>^�j>t�=m�=�        >���        >כE>��p<V׀>y��>��    <1c�=�c�> j?��>�}�>��Q    >ˌr=���        =���=G�1>��l>���                                                                                                L       parents[$l#L       ?���                                                           	   	   
   
                                                                                                     #   #   $   $   %   %   &   &L       right_children[$l#L       ?               
                        ��������   ��������          "   $   &����   (   *   ,   .   0   2����   4   6��������   8   :   <   >������������������������������������������������������������������������������������������������L       split_conditions[$d#L       ?>]R?|�G>����`���j�*�v>Vu���r���ƾ��!�N<f��b�.�Ӽ���=��r�hi=�K]�$�M?z�1i�8օ��y2�����釾�$>�Ӭ�фr�%g~�Wpr>=�r=�,0�O�	>��,�
B�F?w7�@��*��i�j=Kc�;�k�ř*��'=?c8�~��<	{�=����9���Hm;J���Ҽ㴀=��A����8�	J<��@=�蝽%��<�GԻ'����_=�=m�k�L       split_indices[$l#L       ?                                                                                                                                                                                                                                        L       
split_type[$U#L       ?                                                               L       sum_hessian[$d#L       ?C�3�C��aAF�tC��B'%�A$v}@	��C0C')A��"A�`�@]1�@�T.?��|?�B=C��@�?�iiC&JAm^h@�r@�ǯA��?��Y@�l@�^@��BB�|B��C#�\@{XA!@���?�vR?�H�@���@7՘A4չ@��?��I?���@f(?��^?��{?�7�Bc�A)
�?�/�Bѧ�C
�~A�N�@�\F@!�@ml�?��%?���@1�]?�2@?�x�A�5@3�@�|�?�H�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       63L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       %;kh;��
�3�8*�[=���<���n=8>��s&��Z�b=��*��j����=��J>�#�v�> D;����_i>��=��>Է���2>����xU���>f*��)�M��ɑ=��>��3>��n����y�>d����='��L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       %                   L       idI �L       left_children[$l#L       %      ����         	               ����   ������������                  !   #��������������������������������������������������������L       loss_changes[$d#L       %=���=�ܬ    >c4>�gf>>k�>@4�=�H>���>�L>�<4    >Cmb            =�c�=��<�W@=Y@>��=���>"M^                                                        L       parents[$l#L       %���                                                     	   	   
   
                                                L       right_children[$l#L       %      ����         
               ����   ������������                   "   $��������������������������������������������������������L       split_conditions[$d#L       %?�VF?�p�V�i�k�<?;\¾�Q��:M�wK=�Na������������ϻ<�m�=�÷��&�?oM����?@1½�B>՛�>\>�`=�nO���͸�n�=���Klý���<�Ӑ=㢤="����;ͻ��^=����<Is/L       split_indices[$l#L       %                                                                                                                                  L       
split_type[$U#L       %                                     L       sum_hessian[$d#L       %C	��Cƛ?���C :�A�B�PA�W�@fw@�D�B�ahA���@�hA�~�?��?�=@"ҝ@��B��c@�@i|A[�;@p�GA�jx?��#?��WB��`?���?�d7?�]?�N@yu@���@�.�?�#W@$�A]��A8ML       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       37L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       1�������D=Dõ�NJy�7�\�y�R>1ڙ������>�����ʽ��O>
�>�CR=Y�d>�]������77ʑ�:�Kv��W>��7�Z�6>q���AF=�̾X>c����/B=�����6W���w�+O<�]�ͩb=ţj�$�z��>�xk�&D���>�2��L6��Jz9��
���>$���gR� �<L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       1                         L       idI �L       left_children[$l#L       1               	      ��������            ����   ��������            ����   !����   #   %   '   )   +   -������������������������   /������������������������������������������������L       loss_changes[$d#L       1=�@[>P�{>q,6=q�8>b�v>1	�>".�        =�G�>8">Vd>&z�    >4�        >�S>�q�>��5=�]�    <kĞ    =���>�
$>�h7?�r? ��>~�                        <��0                                                L       parents[$l#L       1���                                               	   	   
   
                                                                                       $   $L       right_children[$l#L       1               
      ��������            ����   ��������             ����   "����   $   &   (   *   ,   .������������������������   0������������������������������������������������L       split_conditions[$d#L       1?��\�g�=�G�>��P�a�b��LƾQ⠽���0d�>AA�`���W�@S�=��?�C�=�=2����=����]t =?���=��?��{=�-?�S�<J(�?#"*�* �[��5s����Ͻ�3\�M�;�|p���C<�*�?ܭ��6{�=����G����=�<�u���&,8�8s�.�R=E�������j�L       split_indices[$l#L       1                                                                                                                                                                                L       
split_type[$U#L       1                                                 L       sum_hessian[$d#L       1C��C�Z.A�Yt@�F|C�9A�8AB�@$?���@݄C�YAkN@�D=@P[e@�W�?�&�?��A_�iC��A7~i@O>�@�M@�-?��*@���@�b�A{@ɓ;C��A#�l?���?��?�u[?�ߥ?���?�c�@#?��@$��@���@�g|@��U?�˗@�>RC���@J�@�R�?�2?�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       49L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       /���F;�L��B�~9�h>]Շ�o �|ؒ;CZ��_��>���vv>�R�a��z^<~�辈{����=�b������]�;>�*>��~f�=�;�;o�h���M>am��b�����>���=Mp�~�=>��ʽ��M:���>���>��6�1�x�&� >������n>@v��D���m�:�N>�Q�>S�9�}!L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       /                        L       idI �L       left_children[$l#L       /               	               ������������   ����      ������������            !����   #   %��������   '   )   +   -��������������������������������������������������������L       loss_changes[$d#L       /=�h>�$h>24�>Y�u>*�f=��>WV�>u�<P20<�            >Dv    ?Gw�>�/n            >`��>�X?r >��b    >�?E>���        >R&�=́>,5>��                                                        L       parents[$l#L       /���                                                           	   	                                                                                L       right_children[$l#L       /               
               ������������   ����      ������������             "����   $   &��������   (   *   ,   .��������������������������������������������������������L       split_conditions[$d#L       /?΄?� ?��?��=�G?�J��'k[?iF���?�������}*�����$q��ǰ?a��=E ���� ���=�2z?ʿ&�%V�C14?`BH�.���~�*��Š=�g��1R@�(�%��?��z9ݿ*=�k=��t�Ub��HU�=��O���Q=fw���R_��P�:�b>ʲ=~���{L       split_indices[$l#L       /                                                                                                                                                                         L       
split_type[$U#L       /                                               L       sum_hessian[$d#L       /C���C�}�A�bwC��@�0F@TaA���C�&*@Yt�@~�?��s?�W�?���A�*H?�x.C���Af�1@�(?�qT?Ǚ�@O�AT
A$JvC��M@M�@�u�@�q?�Fa?�Y�A��@��@���@�@C�C�?�V�@�\�?�e�@��F?��@�M�@��N?�t�@=��?�y�@aFZ?֞(@v�lL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       47L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       %;{�k�}�=��:����l��=ؕ���S߻�P�>pD�>4�0<�h�>Q�<���;w�� 9:��>��Ͻ6t�>7�\�ꙴ>1��>3ƾ@�>!#��~>�U�=�}X>���	��<вC��&�>�����p侄Tn�4@���zn=��>L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       %                   L       idI �L       left_children[$l#L       %            ����   	      ����      ��������               ����      ����   !��������������������   #��������������������������������L       loss_changes[$d#L       %=�g�>��=��>!x�    =���=��=�)�    =���=��G        =܅9> ��=�1�=�pT=�˕    =�x�=��-    =gs                     >
��                                L       parents[$l#L       %���                                               	   	   
   
                                                      L       right_children[$l#L       %            ����   
      ����      ��������               ����       ����   "��������������������   $��������������������������������L       split_conditions[$d#L       %?茢?�?J*?��ڽ��@{T?��?Ԑ�=�)F?�-�@M� �dbD;��@?��x�����ɋ@Ij���=\�	� i>���=3
�?z٪=A^c�+��>3q<�0='�J?���;�o����=����TE��˸�XM���_�<��~L       split_indices[$l#L       %                                                                                                                                       L       
split_type[$U#L       %                                     L       sum_hessian[$d#L       %C��B��hA^B��?��A<
�@
߲B���?�~@�K@��`?�\�?�b�Bᆯ@Ճv@�x@B�@���?Í�B�JG@'��?�N�@�o�?�_o?���?���?�Mt?��U@T[�Bad4BW0[?�rG?���@P�E@?Y?ޢ7?�8L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       37L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       E��M'�J��;oq8�!�w=v..�S};���Q8J=@��>*����)��}k�=��5K�<�44�r��=�<����>�>�WQ��6u���`;}���_�����(<L���>]<P:Y>d@���������� >�=�=�
�iO�[$�=��[>����R�Tr�<�r��A��=T/ >���<V�s��ʽ�gQ��W2=��|=�<;>��1>�Pݽ"Բ>�s����q��g=�~���:4�D�=��,>H�K<����Gg��>+�q>��y=*���Gy>�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       E                                   L       idI �L       left_children[$l#L       E               	                     ����         ������������      !����   #��������   %   '   )   +   -   /����   1������������   3   5   7   9   ;   =   ?   A   C������������������������������������������������������������������������������������������������L       loss_changes[$d#L       E=�v`>ō0=ʨ>'�F>��'=�=�7.>��<� >�Vg>7�<�(h    >�`A>���=�$X            >^�>    >DQ        >��>��>���>�&=`>b{<    =�"             =�0h?�4>�4e>��x>��?=�?/�=�̨=��R                                                                                                L       parents[$l#L       E���                                                           	   	   
   
                                                                                         $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,L       right_children[$l#L       E               
                     ����         ������������       "����   $��������   &   (   *   ,   .   0����   2������������   4   6   8   :   <   >   @   B   D������������������������������������������������������������������������������������������������L       split_conditions[$d#L       E� 5D?^�9��n?�a*?���=�5����?��ļ��JA?�S仧I,<=OO��5�?��>�G�<�����=��C!�?����&t�q!��<̽�f0��.?v�>{Dn�$�r?�K����ӭ��P"=dӽ��c��|�?�����@��U>�2˾�
�>�kٿ�/?�$>�j��H��������<���<���=���=�-ּCe�>b��9U�0S�<��ν��r�k����=p�[;�ҽ����*=M��=�+<L
̽��='�dL       split_indices[$l#L       E                                                                                                                                                                                                                                                      L       
split_type[$U#L       E                                                                     L       sum_hessian[$d#L       EC�'�A�e�C��`AsHAw�x@��HC���AFA@3mA�e@��'@��?��C$�C8hA2��?�@�?��8?��@ʽ�@)�|?�K@��_?�5�?���C�.A�ÄC �+@�'�@�i@���?�Ņ@��*?��M?���?�,�@u\gA,�nB�A� �A5�.BJ�EB��@���@�|@�h�?� �@Qt�@6�?���@h�g?��@�@���@��SB���B�&A�@�V@ؐ@�zCB�JA<K�BP��A�T�@oc�?�o?��?��hL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       69L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       ;��@<������N;ة|>��]��:�a <ӎ
��/�=��0?wF>Ҿ�j>~p���M�<��>�X,����=�p���r�>�
��D2��ͽ�D(>�a��;)$�<Ç����Ⱦ	�v��h�=��Z��O���*�=��0��%M>H+T>�Yi�L��	�����>�轺�a���}> "o��T�>]�����C�	����)>L�s>�a�>&�Y>K���R�ʰ����t��آ;RIL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       ;                              L       idI �L       left_children[$l#L       ;               	            ��������               ����   ������������      !   #   %   '   )   +������������   -����   /   1��������   3����   5   7����   9����������������������������������������������������������������L       loss_changes[$d#L       ;=��<?
u�>��5>��>��>��??��>�Yi>p�N        >?�m>�	>�Dh>���>�.;    :��             >��l?C��>t�>t��>��>�P
>n�             >�`�    >ZP=G$�        ;�     >��=X�    >�]                                                                L       parents[$l#L       ;���                                                                                                                                               !   !   "   "   %   %   '   '   (   (   *   *L       right_children[$l#L       ;               
            ��������               ����   ������������       "   $   &   (   *   ,������������   .����   0   2��������   4����   6   8����   :����������������������������������������������������������������L       split_conditions[$d#L       ;�1$��2�b�)G�6�,�z�`�#�'Sп7��?�*G<�f:>![� ]j>�Z�Jy
�!��8^]=��5>i�<�����;=�@[���V?�޿(��?�f?�0�!bԿ=Ʋ��X��%L(���[����Y>�q?�5��_�=p3��(R��u���&�:>���=���ѕ����=@)S����=�N���$j��oe=uċ>:�=Hk=t7��E���:M��~%���:|#%L       split_indices[$l#L       ;                                                                                                                                                                                                                  L       
split_type[$U#L       ;                                                           L       sum_hessian[$d#L       ;C��RB��C��OB���@Y(8A�e�C�4�B�C\@v��?�v?�A�@MF6A��1@��OC�6fBx��?��@5�U?��?���@�eA-m�Aq@�0@��7A��Cy�wBr�)?�O?��^?�qL@�t�@:΢@�� @_-�?��4?��,@���?��?AbLq@���@�tCw�yBJ�3A��?�`�@�\m?��]@��	@=�?��Z@]w�?�Χ@p�VA&@XH�?�5�@X��Ct%�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       59L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       9;�]��Y�=�=�����<���>���TO>�H�%˼;��="�����=�8>y��=�w�/�='��>�����A����<�1;�v�O<�aO>����_��|�`>�|��%�b��>����vC_=*ž(��=,�?���^=}΋����4L�=�U�>Z��͙�=��,r�>q|�<é�������
>~�����^>J���8���=�~����>D�JL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       9                             L       idI �L       left_children[$l#L       9               	                           ����      ����������������   !   #   %����   '����   )����   +����������������   -   /   1   3   5����   7����������������������������������������������������������������L       loss_changes[$d#L       9=���=�i=��p>W�>�n�=��=r�=�*j=;�P=���>�>S�=��=�R�    ><�=�4                =� >�>U    >�K    =    =���                >	'>t�>�?>z &>2z`    =��                                                                L       parents[$l#L       9���                                                           	   	   
   
                                                                     "   "   #   #   $   $   %   %   &   &   (   (L       right_children[$l#L       9               
                           ����       ����������������   "   $   &����   (����   *����   ,����������������   .   0   2   4   6����   8����������������������������������������������������������������L       split_conditions[$d#L       9�%Ʉ�w�h?�t�
nh�f�K?,��>�b��K���͡�� �P7?2R>gEN>,=���b.���<I"N=�ba���u�?����%H=צJ�fX=��e?�hĽ���@.~����nhd=�����<L �J�c�jl��1�><�?�*:?q�n�X[�?Wb=����M<�#�N�==��v;��z��`����=��S��\=�<��sw�2��<�d���W=l&L       split_indices[$l#L       9                                                                                                                                                                                                              L       
split_type[$U#L       9                                                         L       sum_hessian[$d#L       9C��B�!�BB��A.�#B�E�B-Z�@�0�A �@;$�@JY�B��B�)@ͫ�@Y_?�@�ʐ@>�}?��6?��?�:}?�yB ��B0yBA�?�m�@��?��2@�]?��@re}?�_G?�(?�d�?B?IA�A�V	A��;A3�|@ ��@Q2�?��k?�O?�`@�M@zeB�@f�?@�� ?��NA�yA�*@�pv@��G@T�b?��j@�ML       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       57L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       ?���;�j��.)��i"=���=�rZ���r<��B���I���>!�S�}�>��Ͼ���������<�3���Ig<��o��x==��¾S�>K�پ]�J=��=�K�>������{;�$�Q�@�^kS>�<4�¾�_!�ܱ���q=��W=��>�j0>jCٽ�y���Ҽ�V�<v	�O��?�>�����W=f۟���f���O8m>�X=<��̾L�>��S=��a���>^���ŕ>%i�Z�~��L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       ?                                L       idI �L       left_children[$l#L       ?               	                              ����      !   #������������   %����   '��������   )��������   +   -   /   1   3   5   7   9��������������������   ;   =������������������������������������������������������������������������L       loss_changes[$d#L       ?=��{>�F>�mQ=�>��->U&>��$>�]�>�ݒ>��>n�>;W�;妀=��=��R    >E;�?E�@>��;            >3��    =�y        =陠        =���?kw�>eͮ=���>�i?�3?�>4ۂ                    >K��=�P�                                                                        L       parents[$l#L       ?���                                                           	   	   
   
                                                                                   !   !   "   "   #   #   $   $   %   %   +   +   ,   ,L       right_children[$l#L       ?               
                              ����       "   $������������   &����   (��������   *��������   ,   .   0   2   4   6   8   :��������������������   <   >������������������������������������������������������������������������L       split_conditions[$d#L       ?>Dzο����;�>	���X���0��RV�a�Ƚ�7=�I�C�Z��r?��2>�)��/DԽ����i�\>�� ��/����=\��=�>�н� �?�<��=ݍ�?N��:��"�{̴?�t>�06��4L?q�@=4�AG�$�2%]=�m=����_%�����4�?��?�^���=�In�+�<��ƽ�_H�;��x�=��J;���uz�>x2<���3©=����?��==�~�2����`L       split_indices[$l#L       ?                                                                                                                                                                                                                                    L       
split_type[$U#L       ?                                                               L       sum_hessian[$d#L       ?C���C��NB2\WC�8A�q^@�іBb$B��C�@���Ala@�W@$�@�LA�q(?���B�B"3PB�*f@ ��?��?��(AU�\?�ܜ@M��?��?���@�2�?�f@?�IHA�|�A3BӪ�A ��A��B�B �A��@o&,?��?���@o�?�݇AĮ�@�6�@�A�lBR�BT��@�n�@4�0A��?��BJX
AW�@�A�l
@��J@�XA��@��@*�@\_L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       63L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       1�N)[;7Vｐ��:���>�.b�q�/<���<���/����������.=�0:L%�>�DJ�V+I�ӌ/=�׾xH�=Q徢X�>}j?�JW�<kj;�J�W�[
>�+�=iX����>�]ü\F�>�	�=5��Z�=���E.=nԆ�f���0�=ϐ㾯b�?�N>9y��H����������=����doL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       1                         L       idI �L       left_children[$l#L       1            ����   	         ����                     ����������������      !   #   %   '   )����   +����   -��������   /������������������������������������������������������������L       loss_changes[$d#L       1=���>> >�c=�|�    <�,>�(?$�>9�y    =��L>1>3�>���?>�y=�� ?"�                =sd�=�Jm=���>͆>S��=�@    <�<�    >�A        >�t                                                            L       parents[$l#L       1���                                                     
   
                                                                                       !   !L       right_children[$l#L       1            ����   
         ����                     ����������������       "   $   &   (   *����   ,����   .��������   0������������������������������������������������������������L       split_conditions[$d#L       1@�@
�1@,-��W=�7�@"��)��%J��3O���|�@'�>�:k�?�{��.婿)c�	���-��=ׁ����<z���Ъ@<�@SR�>.���fR�4��?s�D<8���> ��.=��?<<�Կ
=�;�)�8<�LQ�0ᓽ�p<�D��v=>�=!Ž��˕󽷰���J_<�#���ERL       split_indices[$l#L       1                                                                                                                                                                                   L       
split_type[$U#L       1                                                 L       sum_hessian[$d#L       1C��sC���A`�UC�@�?�v@�@�A�C	�OCV�V@$rC@
�@8U�@ͻ9C"�A
;@`��CS7�?��?�/?��&?�$c@J�F@P�,B�~0@�p�@"��@�#?�B�@H{@��CP�?�M?�@@��?��B��5B%+�@3G,@��Q?��W?��x@��&?Ꮺ?�yc?��@��QCL�?�,?��SL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       49L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       ';_gw�rw==D��nZ��{>?#�<�-<D������5��>��H>e�Z;���'>@ݾ3��=@���p0�<�M;��ƾs]�>�q=��L�r��=D��>)Pg��m-�N��=����y>&뾖i�=<�w�(�=�/Ǿ�\�;���>%N�<�7@L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       '                    L       idI �L       left_children[$l#L       '            ����   	         ������������               ����      ������������   ��������   !   #   %����������������������������������������L       loss_changes[$d#L       '=�3�>�~=�vP=���    =��=��>��>�j            >
Wx=�(1<�p>�x=:ؤ    >�=�ֈ            =���        =��q>�V!=��                                        L       parents[$l#L       '���                                                                                                                    L       right_children[$l#L       '            ����   
         ������������               ����      ������������    ��������   "   $   &����������������������������������������L       split_conditions[$d#L       '>:	=��I��=�Vѽ�����>{a�?�V?�]׼Z5=�$=��j>��a?2�<�v�@�~�o�T��W���r�4���(=��<�e�@��<lw=K-I?>��??���)8�=)a罴~�<bH)�Jt%<�#��o:��M=F^k;�BML       split_indices[$l#L       '                                                                                                                                                L       
split_type[$U#L       '                                       L       sum_hessian[$d#L       'C�$B��sBI��B��?ô�@[vB<3B�I�A=5�?�V�@[�?˶VB5��B���@O�@�;@�ީ?���B0ÔB���?���?��@ @���?���?��x@SMA���A��PBr�@�z�@�_�?���?��D@�s@$�Av�@��A�n�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       39L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       '��v�<	^������m�>�;���$����;��Q��>�?��`%��
�=Ɯu���q<q7�d��>�m��e/>��?.��>-�>�JԼH��;�(
�:|
>ŉ�=�)��u>:�o�6�< Ro=�~t��e���
>��S�3�s<�>���=��TL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       '                    L       idI L       left_children[$l#L       '               	               ����������������      ��������������������            ����   !   #   %����������������������������������������L       loss_changes[$d#L       '=�h�?j��?O�E>߰c?`b\>⇚>��?+uU?:��=��                ?��>v/}                    >
7>��>?I�?�I    >2	>ӆZ=�                                        L       parents[$l#L       '���                                                           	   	                                                      L       right_children[$l#L       '               
               ����������������      ��������������������             ����   "   $   &����������������������������������������L       split_conditions[$d#L       '�3���u��i��&�>�%<�ٔ��������n=�c
��|��&iA<�UZ���=nO��0�2>A��(yl=>�->Q�=P�|>�/�?�ҿYR�?��=����xN����>�|�[bl;@b�<�1X��ɽ-h�=��1�W֋; �$=�)+<���L       split_indices[$l#L       '                                                                                                                                                 L       
split_type[$U#L       '                                       L       sum_hessian[$d#L       'C�j�CgB�B�%
Cbs�@���@�	�B�$qC]��@�e�@g��?��]@Z��?�4�@Y��B�X#C\9�?�y�@(/�?�8B@'k�?���@�5zB�d�CV$@ºQ@}�@!b-B��@�d@��VCQ��@f
F@j\?�l;?�XAl�xBW�?���@�2�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       39L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       ����;�V���=�!�9��	�#��=�o��d>��e�F�;C5��&΁�g�t���Z�;Q�K��q�>Tw������B=��+�nԵ�����j%G>�oh�v��;&}о�����;=�����L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L                       L       idIL       left_children[$l#L                      	   ����   ����            ����������������      ������������������������      ����������������L       loss_changes[$d#L       =�[z=���=��r>j��>;3�=&�T    ;�%�    =�;�>`�;=��z<�0p                >)_�>`�                        <��=�Q                L       parents[$l#L       ���                                               	   	   
   
                                    L       right_children[$l#L                      
   ����   ����            ����������������      ������������������������      ����������������L       split_conditions[$d#L       ?
ڿo�|>����p���m����X<ƅU��p�=��࿂�j��?o����=8�ý��5�:{ˎ���M�|���it5�66�= @���Lm��ּ�|�=����6��`ن��}����<�2����L       split_indices[$l#L                                                                                                                           L       
split_type[$U#L                                      L       sum_hessian[$d#L       C�%�C���@��7@���C�$�@��"?��Q@	b@A��@sa�C�=�@U@4��?���?��?��]@"��@�I5C�(�?���?�<�?��A?��?��,@4��@/ZWC��?�a�?�S!A�w�C��L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       31L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       3;5��� %�=ML!���(�D�>W�<]}�0D=�**��澁:�;��9>��=d���ks�<����)>"���=�X=����z�%Ƹ��T�;�CK>N6*��\�<���>��L����A�"=�:�<��>L���Jۜ=Z�\<`_+�,�u��fA>�.��9��yy޾	��>F�> ��>��`�<�=��=����>��<��	L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       3                          L       idIL       left_children[$l#L       3               	            ����������������                        !��������   #   %   '   )   +   -��������   /   1������������������������������������������������������������������������L       loss_changes[$d#L       3=�(M>MT>m\=���<�`�=�8h>k`�>�=�?                =�
=��>��=� >&�8=�M/=��H=��<        =�2=�$�>6��>8��;�@=U��        >Rm�=G�H                                                                        L       parents[$l#L       3���                                                                                                                                                          L       right_children[$l#L       3               
            ����������������                         "��������   $   &   (   *   ,   .��������   0   2������������������������������������������������������������������������L       split_conditions[$d#L       3?�7�?��t?�t?����s.>���?dk���?�0ʼ���h:��=�0@,�?��&?K�>��>G�H?�@J���+�F�w�ǘ�>�\=_���Z�\�%?�Ɓ?o?|�h��=��?өǽ&�T�sm�<�L�;����O;Z���=�k�^[�����%f�=�=Ǝ=�$t�0�0<�V�=p��7Fk=��q;��L       split_indices[$l#L       3                                                                                                                                                                                            L       
split_type[$U#L       3                                                   L       sum_hessian[$d#L       3C�UB�E�A��BԦ@3��@`��A��B�o=A�:?���?�2?��@A�@'�B�x�A���@��@F��AhO,@O#�?�O?�8B~Oo@*"A��A�{@eqV@x�?��J?��AѨ@��?��X?��[Bus�@��?�&�?�wA�@�@�ܪ@N��@�(�@	�)?�Y?�_�?���@���@e�&@fף?�<�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       51L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       =�3�8���t<
̜�Si��M�;��>�� �AF1>:�5>i�輼�U�4@=/���e��=S�=$(�>�q潷=E�<�Fý�(�>*��<Hg�����;ʔ�>9�q�w\�D��=@�>ٴ$;��>?�;�d���;�o$��aD>o뼟��>U;��l���-��p\�B�_>2��(�=��J��
�>�@C�'��>k���>��S�!I���l>�h�>��A>!l=Z/*�U�dg>��L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       =                               L       idIL       left_children[$l#L       =               	   ����   ����               ����   ����            !   #   %   '������������   )   +����   -   /   1   3   5����   7   9   ;����������������������������������������������������������������������������������������L       loss_changes[$d#L       ==��p>��s>5D>g>>��x>
ܙ    >�0    >�h>p��>��">�Y|=�g�    =��X    >�[&>؆�>�e�>��e?Z�>�x�=�K�            >��4>ӟ�    >U��?5>�,">�ن?QY�    >t��?B>/}.                                                                                        L       parents[$l#L       =���                                               	   	   
   
                                                                                                     !   !   "   "   $   $   %   %   &   &L       right_children[$l#L       =               
   ����   ����               ����   ����             "   $   &   (������������   *   ,����   .   0   2   4   6����   8   :   <����������������������������������������������������������������������������������������L       split_conditions[$d#L       =>�]9�U�*@��@<_�=e2�>�7l=�'Z?�R=`W=F��=3k����^?)��?��<~��T��=ꈮ��_�=��@�`
�����y��.z�H�,:��=^ꈽ(�<?=�m?�r>�I���>���?D��f�l>h$z��R�[K��?*t��*����j���	�i�=V~�J��<��Y���t=�淽I"y=����=���AC%���O=���>'�=��<���>�ͼ��q=���L       split_indices[$l#L       =                                                                                                                                                                                                                           L       
split_type[$U#L       =                                                             L       sum_hessian[$d#L       =C��1B��`Cr��A[�Bz��CqYe?�&�AK 0?�\z@���Bh5C,/"B�T�A1�#?�xe@)	?�A^A��WA�B��B�G`AM�BaHJA��?��?�lS?���Aft�AK�?��AꎪA��B��B�OA�\�?�`A4!ZBD�@�@ؼ�@!qM@��^@���@�8&@���A�]�A:a�@�p�@-&�@���B�F�?��KA���A�ۛ@�%@H]�A	�B��A�AE?�G�@��L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       61L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       !��լ:�%q��,Q;BqW��Q��ɻ�|D;�-o�,rѽZ�0�5�ĲC=�'%;E�	>W�i��;Q���(;��d�@�D>��ƽ|�_���#=��;>�}>�콅l����$>�H�=�W5=E�u�H�>>����$L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       !                 L       idIL       left_children[$l#L       !               	   ����      ����������������         ����         ����      ����������������������������������������L       loss_changes[$d#L       !=�U�=��'=�5H=}p�;��0=JS    >��>]�                >��>ֆ>�g�    =��<��8<��    >�С>�ZL                                        L       parents[$l#L       !���                                                                                                  L       right_children[$l#L       !               
   ����      ����������������         ����         ����       ����������������������������������������L       split_conditions[$d#L       !?�	?��R>�� ?΄���i��M���\?��=�[�0҅�S�s��	<�ȓ?��L=�C���[��Ɨ?��M>�ŵ�Ve����?��r�L,W:d�0="�������$�=劝=g�<m&�p��=�������L       split_indices[$l#L       !                                                                                                                      L       
split_type[$U#L       !                                 L       sum_hessian[$d#L       !C�HC�f�@��ZC�A�@��@]��?�-�C���A؟<?�JY?��?�i?�HYC�9e@��A�
t?�L{C��@E��@sc�?�`qA�?A�kC�j@�hB@W�?��y?߽U@�-@�SA�@�
�@���L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       33L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       G;�R���=K&�<z�]�J�>C��<҂ɻ�-�=��%�7J���9>�<�T���?�=��a<?a��(>�J<=_f�'_�=;�>������=e�Ѿ�>=(
���d����>L�N���H=���;���>;�h��Ǿ=�ھYaf���j>Q��&�ʾi�=��>�S<�N'=���#/W�u�9<���>�Q�<�ѐ���5����=�"�^��>��r�-��C�>	�O�ar�= {^����=!챼m��>��<�1�]}���
:�k� �H��=���>o���I��L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       G                                    L       idIL       left_children[$l#L       G               	                  ��������            ����      !��������   #   %   '   )   +   -   /   1����   3   5   7   9����   ;   =   ?   A��������   C   E������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       G=��g=�O=��=�>.N/<��p=��=�T�=��=e� >44%        >%-�=��F>�>'�    =�<ٟ         =�{y>��>,�=�w�=݈�=��y=P��<I�@    >J�A=��=�R�=�28    =���=�ΰ=��.=j�        <���=��                                                                                                            L       parents[$l#L       G���                                                           	   	   
   
                                                                                                     !   !   "   "   $   $   %   %   &   &   '   '   *   *   +   +L       right_children[$l#L       G               
                  ��������            ����       "��������   $   &   (   *   ,   .   0   2����   4   6   8   :����   <   >   @   B��������   D   F������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       G?GĿd����:�zH=��E>AA�?��2������:@��>�=�;똤?��?�+?[/D�� g=�Y�y��"�<`j�=�I���e�R:b@*�>���?���2)|?���U_�<Ù�Q?�*u�-���鬽�m�?�K�����>�t�P��<�
=���?�[�?p,0�C�i��r�;�s^=���;��z����Ŕ�<�4�����=��V�P�t�k=%i���D�<-���N�<BO;����=ï1</뽄�������] �p��<���=��ʼr*L       split_indices[$l#L       G                                                                                                                                                                                                                                                               L       
split_type[$U#L       G                                                                       L       sum_hessian[$d#L       GC^�B�&8A�]�B��B vQ@ 7A�]!BL��A}T�A@��A���?���?��A`��@��SB9�x@�c�?�Q�Alj�A0v�?�'�?�>&A���A�@���@�T_@m=�B/��@\�@A+?�7�A7��@R�9@/�A��?�oA��\@Kg�@��M@r��?�V1?�� @>/@�4?��gAn#�A��[?��l?��.?��W?�o�A{@�@�-?��?�t�?��J@���?���A"s�Aq_$?��?���@�j�?�6'?�E�?��?�s�?��?�:�?�U�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       71L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       7:2al��R<��ֻ4���d~!>r?;�̻��>�]�=�����,�>b'ʾe��M�<ܹ���S�8��o����;��b>�M?���>;ؾ��;��>��<,q�DH�=��$�a��<D�n��O�=��,>�¾| l=R)�>�k��� ��>��л�F��r��=�(�>ى���ɻ�D����A>�:�;�K�>�Ye�1�}�����O��<�n�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       7                            L       idIL       left_children[$l#L       7               	         ��������                        ����   !   #��������   %��������   '   )   +   -   /��������   1������������   3��������   5��������������������������������������������������������L       loss_changes[$d#L       7=�,N>�/�>P�K>�s6>|�,>�O�>�Q>5�%        =��P>��F>��=�J>�Z�>@> -c>Y�    >h�=�Px        =�_x        >��4=��<<��m?�b>���        =��W            95�         >�l�                                                        L       parents[$l#L       7���                                                     
   
                                                                                             !   !   %   %   (   (L       right_children[$l#L       7               
         ��������                         ����   "   $��������   &��������   (   *   ,   .   0��������   2������������   4��������   6��������������������������������������������������������L       split_conditions[$d#L       7?0\�?#�@�W4�?П>AA�?c�̾����=�p�<�E�>�t��%�?��ҿ*A+���?�a*�&���-�ʾM作3z����}�=`��=�k:��^=�?9�?��ľ���(�ѿ%�G���R<�F5?�&��F�<|2	>���V6�O�=��<��Ƚ���<���=�e�\a�Ɂ�=��T:��l=�ѭ�U[ʽ!�|����yhU;��(L       split_indices[$l#L       7                                                                                                                                                                                                  L       
split_type[$U#L       7                                                       L       sum_hessian[$d#L       7C��Co�*B� &Cj��@��tA>�B�O�Chě?��?��@`JmA�r@b�@���Bk(�A!�C^��@"C?�PT@���@��??���?���@���?���?�"Bcϗ@��@��B'�sC4�~?��>?��G@1�?��+?��@�2@4�?�g?��B^*@Ԑ�?�k?�f�?�?ABڅ@�Om?���C3?�?б-?� @?��^?�8�@�
BI��L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       55L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       =��<����<.]t>�w{�����t<��c����=�O]>��>�����>^�'����=��C�h���h>���2�K��h>��<㼇��391�=Nצ�4��m=��[=��V���e�޽�=��>O�ɾ�噼��ؾ���=�YǼ.Wռ���=̓h���=�����>:�3��Ҿ�����^�����+>��>�e��w<�>>o������ཌ�>
Lf�� ���Kz��!�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       =                               L       idIL       left_children[$l#L       =               	         ������������                  ��������      ����   !   #   %   '   )��������   +   -   /   1   3����   5   7   9   ;����������������������������������������������������������������������������������������L       loss_changes[$d#L       ==�>Δ>r&�>���=�E�>~Æ>��>K_�            >u�>Q��>{�L>X��>8j�>�        >�j�?"5Z    >�">��>��a>Q�>O�?        >���;��=�i�=,��>;�     >�|�=~>���>�Ǵ                                                                                        L       parents[$l#L       =���                                                                                                                                                             !   !   #   #   $   $   %   %   &   &L       right_children[$l#L       =               
         ������������                  ��������       ����   "   $   &   (   *��������   ,   .   0   2   4����   6   8   :   <����������������������������������������������������������������������������������������L       split_conditions[$d#L       =�1$��2�b�)_�4D�,�z�`�#�'Sп�s��jf<��p>D� ]j>�Z�I y�!��@|?.P���=�A����V?��=�*�>�Ӭ?�0�z�]��?��J��p�<��n�[��g��>�q>2� ?�{���F��UB>���@����Y����<�����u�=B��Ŝ=`>�rK��놼�>����+z�=:��=��^��W�=d�	����a���=%�H���н��-��(�L       split_indices[$l#L       =                                                                                                                                                                                                                             L       
split_type[$U#L       =                                                             L       sum_hessian[$d#L       =C���B�(C�-�B�i@S�A�7
C�gB�4�?ң�?�_*?�Э@B�A�ؓ@��FC�C�Bt2�@Cnt?��p?�bA"��A��@k�j@w#A�B�Cr��Bi!�@1�?�Y�?��X@���@.*@�#N@Z��@/��?��wA[q?@�(�A��C[��A�EB�"?ߞ�?��@?���@���?�I�?�
P?��@�jl?�=.?���?�AQ?��~@�̣A
�@H�g?���A�u�?��	?��CZ L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       61L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       1;EV����<���?f]����dg#=(,N>f�z�䘻�x�>�I>�8Q=8N�[�-<�ƽ\��>><���Md<�RF�G5�=a��#�^����>_�2��֍����>R��p-~=?U�>\<�8���c����h���>x�>���0I{�ew�=J�����}�a<�����p&=�<>�5u=��>�3�<�=��L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       1                         L       idIL       left_children[$l#L       1         ����      	   ����         ����            ������������            !   #   %   '����   )   +   -   /������������������������������������������������������������������������L       loss_changes[$d#L       1=�ݵ=�׎>62    >�=�qB>��    ={m�>	��=ε�    > @>/�V>��=�{            >�BH>�e�>�>,;�>U�m>/�>�7    =�V�=�dY>P+�=��t                                                                        L       parents[$l#L       1���                                               	   	   
   
                                                                                          L       right_children[$l#L       1         ����      
   ����         ����            ������������             "   $   &   (����   *   ,   .   0������������������������������������������������������������������������L       split_conditions[$d#L       1��8�w��29D�e�
��ʿH�!�-Wz=�|}>ѯ��XCe�d��=�b�c6;�B�/ ��Q��=dHܽ��;��:2�A>ؽ�M�>
+u���I���o�kĨ=/�xt$�Z�Կ"e�/�����ֽ�۱��x=�\	=���S�a���J<s���3�\��.�;�+���Sa<���Y��<�SX=�pn�b��<*2�L       split_indices[$l#L       1                                                                                                                                                                                 L       
split_type[$U#L       1                                                 L       sum_hessian[$d#L       1C��B?gB�K@�3B7
(A��B��(?�e�B16�AH�!@nS�?�=sB�P2B��A5	A)�
?� �@:m?�2�Ab��BI��A�uA��2@l�@�AE?���@��"A�.@�>�B*� @�nY?�
BA�TI?���@��?Ԅ�@J��@�G�@ׄy@>?���@G�vA�n?���@��	@@�:?ↄB#y�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       49L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       E:�� ;���;�:��=�����=N�Һ߽�>$��jY>=0�����>9y<>5 =����:-���`��>W*^��O�%C�>	"�=B�>�M��-�5=35C>kw��u��1�<�^��	�U>9��Ь�>�7x=ޝ���>�`��`^w>!��N�X�}b~�eU�>C�~��G=֞>�|��t&��a��>p�}����:ưG���'>�Y�<s^?>?]��"��.>e&��WiE����=�e)�?�}>��)�5���g��= �>�����_l�3"X=�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       E                                   L       idI	L       left_children[$l#L       E               	                     ����         ����   ����   !   #   %����   '   )   +����   -   /   1   3��������   5������������   7����   9   ;   =   ?����   A������������   C��������������������������������������������������������������������������������L       loss_changes[$d#L       E=�C|=�f>z�4>Ú>��#>5�&>��e>-�=���>L�>��>GAX    >U�=���=�    =���    >�>�=��~>��    >hX>$�1=��    =1/@>$ՠ>�r�=8��        = ��            =彸    >�!>>�!=�^�=�W�    >��            =�[                                                                                L       parents[$l#L       E���                                                           	   	   
   
                                                                                             !   !   %   %   '   '   (   (   )   )   *   *   ,   ,   0   0L       right_children[$l#L       E               
                     ����         ����    ����   "   $   &����   (   *   ,����   .   0   2   4��������   6������������   8����   :   <   >   @����   B������������   D��������������������������������������������������������������������������������L       split_conditions[$d#L       E>Dzο��=ԥ�@
��?'<z?��.>��?�A|�ZJ�>��V�2�J?�j�=^�|?��E?6��?�r������ܻ��x�B�?7Pw��9�=�)�?��?ԼL��D��d?>o�w?�q?؉����T��h�=�uľ��)���9=�@ʻ���D�½x��8p���?�ѵ@*
<04�?P����}���g"=�k�?�4r9�m#���b=�w;�Y=e����D8=�}���?*��`?<���e�0=�x��ZQ���F<��=�Dǹ���V�<>c;L       split_indices[$l#L       E                                                                                                                                                                                                                                                           L       
split_type[$U#L       E                                                                     L       sum_hessian[$d#L       EC�~C�"�B'��C{��A���A�,yA�Cv�@��@���A&T�A�s�?���A��Ad~CuG�?���@ayg?�C�@�Ws@,t�@�-@THA���@��@Բa?��@_��@��Cr�0@. k?��]@ ~8@X�@BU�?�$�?���@� |?���A9��@̰�@�e@$��?�U�@��@	�?��(?���@�.�Cp��?�%?�}�?���?�Gc?�j|?��4@���@p�@��~@�6�?���?�@?���?��]?�X�@}CU?��B@��@d�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       69L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       ���9֨ҽ��b�ܺ<=�-`=6���9e������!.>�"��T?I=�	+=	�&�VUk���>E�P=[n���]>��=Kj�)�ƾ��q:��پ.T�3>-`�=�vP���L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L                      L       idI
L       left_children[$l#L                      	         ����      ������������      ����������������������������      ����������������L       loss_changes[$d#L       =�gJ=�y�=sߦ>S��>̹�<�5=�_�=�V7    =�OY=���            =K�>                            =ɩ�>g�/                L       parents[$l#L       ���                                                     	   	   
   
                        L       right_children[$l#L                      
         ����      ������������      ����������������������������      ����������������L       split_conditions[$d#L       ?�2?�����?��Q?^������?z���y�;���q�%�~�X<�qg<%3Ⱦ�@?IK0=m�a<��i��!�=���<��K�����"?9�ξ�~s�;��=P�<�Zǽ���L       split_indices[$l#L                                                                                                             L       
split_type[$U#L                                    L       sum_hessian[$d#L       C�ۓC��9@�V�C�+@��}@"1@�E�C�}�?���@'>@S��?�m&?��<?Ǹe@�WvC���?���?��?�c[@$?�I�?ٛ�@��C��t@r��C��^@��?��2@WwL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       29L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       :a�&�L��=�:�N�
��E�n>WTy��0=�Mv�R�a��ם�Hf�W�z=��\�$���q�>Q.�>@v�csF<x�ҽ%�>b�:;�	L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L                   L       idIL       left_children[$l#L                      	��������      ��������   ����   ����   ����   ��������������������L       loss_changes[$d#L       =o�i=��=���=���<��h        =ԤR=��        =��J    =��~    =���    =�oj                    L       parents[$l#L       ���                                                                    L       right_children[$l#L                      
��������      ��������   ����   ����   ����   ��������������������L       split_conditions[$d#L       @*It?�����L.?蠦?�pD�m�Q=�2�?�@X�ӽ}1B��W?��ڽ�b>�Ӭ�)_��d�={ǽ��v��x^;�N�F)=��#;�L       split_indices[$l#L                                                                                        L       
split_type[$U#L                              L       sum_hessian[$d#L       B��zB�1@Z	B�?@_�;?��?�0xB�A8Yo?έ�?�N�B�)K?�q�A&Ҕ?�6�B���?̙EA�?ǀB��dB(�@��1@rO�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       23L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       ;:ػ���>�<%<W���9��S;�[�>�cU�LS�=��1>8:C���>AW�;�R��m�<�ր>"�(����>�l@�k�P�#�<%'>��a�7�h�U{F<�����.]���E>�r�<�����3=%D�>���Nݾ�8<�K�>l�;�I	���t����.�.=�'�>$C�������=��>��I�f ���d>�tY�T�=���=�]�e>��ἤB
>���3���^�<�ayL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       ;                              L       idIL       left_children[$l#L       ;               	   ����                     ������������   ����      ��������   !   #   %   '����   )   +   -   /   1   3   5   7   9����������������������������������������������������������������������������������������L       loss_changes[$d#L       ;=��n>Y��>�W>H�D>���>\�    =�\$=&%&>�->�`�=���>2��=x$�            >��    >v�`>�H�        >��9>�հ>X�=���    =ֹ=>6I>l�>��0>4t�>�V�>���=�Hx>�!�                                                                                        L       parents[$l#L       ;���                                                     	   	   
   
                                                                                               !   !   "   "   #   #   $   $L       right_children[$l#L       ;               
   ����                     ������������   ����       ��������   "   $   &   (����   *   ,   .   0   2   4   6   8   :����������������������������������������������������������������������������������������L       split_conditions[$d#L       ;>�]9�U�*@��?�s}=��>�F=�D ?���@-�z�� g>�������,��?�8V;��4=CV��S�<(g����ʾZU.?	�=��B�\4�>�7l�(���w�v�u6�>x<�[�?2g?��>;&龍��R48?^�?�,��&x����1�6�Qqk<���=E�8����U<�H}=�3��<������>	���<�!�<̘׽�t�=�pB��=��¼W�����4;�t�L       split_indices[$l#L       ;                                                                                                                                                                                                                 L       
split_type[$U#L       ;                                                           L       sum_hessian[$d#L       ;C�)oB�uECl�<AO��Br�gCkm�?�MAX@A�@���BX]�@;��ChA	i�?�p�?�?��@�M?���A%8~B/�?���?�SAB,�C=O�@�y�@@��@:��@�>@�$z@l�@6r.B#�sA���A��1A�BC4�1@g�?�k�?��?�а?�sW?�[%@�nT?�ؘ?���@%?���?�>�A��A.q�@���Ah�@�uA��#@�T?���A�^C,�kL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       59L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       =�熟9*8����;����&~��1پery<�+'��t=B���������=�)y;�ʡ>�T۾*\�:ƍ����=�%� h�~ݏ<�-˽y�t>���=X��>'�þ~�t>��8��h='Y���C��$�>V����>���=�D0����:�Ş>,�>H�����2>��p>8>�!N	>��&="%���0��=z>��>�Ƶ���iƼTS�=�N>T���d@>��K;�=^���R�
�����@L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       =                               L       idIL       left_children[$l#L       =               	   ����            ��������                     !   #   %   '   )   +����   -   /   1   3����   5   7   9��������   ;������������������������������������������������������������������������������������������������L       loss_changes[$d#L       ==��=���=ra0=�p�>? �=��    ?��>�E�>2{j>�f^        >�a>���>��3>��=�Gw>~�*>��]>��>QJ>˳~=jTP>�     >�Y�>��>�~�;߂�    >���>A��>�ό        >6I�                                                                                                L       parents[$l#L       =���                                                     	   	   
   
                                                                                                                 !   !   $   $L       right_children[$l#L       =               
   ����            ��������                      "   $   &   (   *   ,����   .   0   2   4����   6   8   :��������   <������������������������������������������������������������������������������������������������L       split_conditions[$d#L       =?�	?|�G>�� �F��8�ھ�M�����&0��X?@1¿H4��㩙<�1�>�� � �f�,��e�� ���L٨>�{X>��==)�?6M?P��=Iq���RB�����V�, ;��"��C�Ӿ� �0Z�=�i0<ڸ:�qn9���='@=q&���>�D=]W�A��=�Ɣ<B����l뺣|�=�c��s����~��<�]�=?2Ľ��=ř':a�<��g�}&��Ӿ��L       split_indices[$l#L       =                                                                                                                                                                                                                                L       
split_type[$U#L       =                                                             L       sum_hessian[$d#L       =C���C�5@��IC��fB&w@U�<?� �B��CC�^Al��A��?���?�X�B���A��A%|�C9��@l��A1eA���@�5PB�QA�f@���@�>�?��A��@a�XC6
M@b�?�q�@{$-@�7�AdI�?�J�?�d�@��B�0�AGvx@|�MA��<@#��@;�8@��@�@<@�+�?���@��?�>,C4��?���?��q@q?�+x@�l�@7��@��@�~�@E�@C�iL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       61L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       7:��=��h�<�w��:���W�P	!=�j=�z��"��<�|���>�H&<�a>�������J�����˽��>Xt��x��>#7A�>�=Ndc�.�>9����I<E�\<��𾄔�=3��>�y`��Ft���I�Xֵ=��>Q3<�}A��C�=[{m�Y:�G�->A��>���#=����������7<����p��h�>>h�=�.G>����3'�=m��L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       7                            L       idIL       left_children[$l#L       7         ����      	               ����   ����   ����            ����   !   #   %����   '   )   +����������������   -   /   1   3   5������������������������������������������������������������������������L       loss_changes[$d#L       7=��=��=�sj    >m�=�sV>8N>�=�h�>r��>ft�    =�.�    =�7k    =�qQ>"�B=[0=sp�    >^>u��=��*    > X">���=�/�                <- =��b=��>-y2=�/�                                                                        L       parents[$l#L       7���                                                     	   	   
   
                                                                                   !   !   "   "   #   #   $   $L       right_children[$l#L       7         ����      
               ����   ����   ����             ����   "   $   &����   (   *   ,����������������   .   0   2   4   6������������������������������������������������������������������������L       split_conditions[$d#L       7��8�w��29D�_GM���ǻGϬ�-Wz�T��G����[�K�n=��ȿc6=��L<E�N�s	K>;w��(h�a�=�kyl=C�辽:2�A>ؿcX=1��0����ٿNv4���<W��=������Y�ʿz�r�sD�"e�1�����4<��u��V��o�=1糼�����=��ج_��+�<	���i�(}�=d}�<��"=⃍�V��<��NL       split_indices[$l#L       7                                                                                                                                                                                                           L       
split_type[$U#L       7                                                       L       sum_hessian[$d#L       7B��"B;��B�ڦ@ �B3��A��	B���@���B�9A*�@��/?��LB}(u@�@O�^?���BQ�@�N<@;�r@�8?�H�A`'JBE�@��?�L�A�`oA�Cs@���@/P?�w�?�'<?��3@J&@��KA�$@�QZB'Tw?��n?�oA3A,@��eA�JAL��@=@S?��?�Kd?��s@LP]@�z8@+� @�0�@*A�A�i�A�?AL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       55L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       E:���	��= Đ���Ծ��[=w�]�!�	�ҦA:^��=��=��w��O�C=K�p<��m�>��C��>�=�G>�q>D3N��!��\ٽ�fR>��S�ȵ>V���#����v9���=��>�T�!��>-�\=݉�L2��g�>������=1x��;B�=���=�V�>���H>x��<��1>��=�m���6|>=��:_ݽ���:ȑ�>����s�=&��>�^l��r�=�%�p(�=cJо�R'<��>cb�& ��N�u�����I�4=��EL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       E                                   L       idIL       left_children[$l#L       E            ����   	                                    !����   #   %����   '   )   +   -   /����   1��������   3   5   7   9   ;����   =   ?   A������������   C����������������������������������������������������������������������������������������������������L       loss_changes[$d#L       E=�K�>r<�> f`>��    >ks�>��M>u+>�c�>��A>�[>Wd>��>�f�>��<v >Y:�>yEv    >�C�>��B    =�RP<�B >`S/=X�>-��    >/!�        >I�>�L>�
D>*�=�e4    >4��>�|�<�V`            >�3�                                                                                                    L       parents[$l#L       E���                                                     	   	   
   
                                                                                                           !   !   "   "   #   #   %   %   &   &   '   '   +   +L       right_children[$l#L       E            ����   
                                     "����   $   &����   (   *   ,   .   0����   2��������   4   6   8   :   <����   >   @   B������������   D����������������������������������������������������������������������������������������������������L       split_conditions[$d#L       E?0\�?.�?��D����n?��ÿL���V�X�@N�?�����?C�X�AE?o�R����>P�?��>w�=�T��o��?ڈ����?
X�0�>�E,>��H����6�?��z<���=��{���?#�@�:�q?$��=5&<=��?���@ ^�:�"<���<�h!=��-?��=�<�;Ыo=���<������=cxt�_�=��X�9��=�*f�0�<G��=�������<��E��l<�`���/;,;:=�n�GZv�xb'��lr�r=-�L       split_indices[$l#L       E                                                                                                                                                                                                                                                      L       
split_type[$U#L       E                                                                     L       sum_hessian[$d#L       EC�r�Ci,�B�qCg�7?��7BQ��A��\AL/�C[,>B	��A���@�AAd@ר�@���@(\CCX��B�@ @�:�AIy�@1�K@��@'�A:�@W'�@X)�@<�4@D��?��?���CR�@���A��x@aH@�m@M�{@� �@���@UY?��?�Z8?���A!��?�ev?�'s@�?��+@Or?&?��A�P�C9�@0��@BݤA�;�@��@	e�?��h?���?���@���?��6@D�@/��?�ȉ?��)@��t@j`�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       69L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       ;���,:�(���_�<[3M��7X=�����9;�ϟ>�d޾��c;�/>^���mCm�m�F<i��=uq��"�>�­=��0�t��ڰO>2o��K۾�Ry��K><����R<v��>�N��v�����C�rv�>��� ⨼���)�H>����V��X㽯�^��i=2�>-�W<�o��+<��\?	o��]>��@>�y����-��������>f�̾���>�
>��<E�W�O�]L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       ;                              L       idIL       left_children[$l#L       ;               	                  ��������            ��������      !   #   %   '����   )����   +   -   /   1   3������������   5   7����   9��������������������������������������������������������������������������������L       loss_changes[$d#L       ;=�)=���=�{�>�d?oz=��$>'>`�>u>�Q*>�)        <�mP=�\?0>�j        >��G>O�>�^t?n�;ث�    ;��x    >V
�>M�l?i.�?��=�<            ?�>2R,    >�8�                                                                                L       parents[$l#L       ;���                                                           	   	   
   
                                                                                             #   #   $   $   &   &L       right_children[$l#L       ;               
                  ��������            ��������       "   $   &   (����   *����   ,   .   0   2   4������������   6   8����   :��������������������������������������������������������������������������������L       split_conditions[$d#L       ;>]R�/�Yq`�=�y�ZH�<lgA��à��z�=�k�,�j=��$=��o��[�?��j=6���������>t�<���?-F�>�f$�UW =�ƿ������>��� 2?@f�Y��=S�����4�VgG=������ě�?K�^�>($� r>�)мҾ�à<4<�=Pr<���>�<<>$볾�=��M>❻��j��+���W�=���״ >
��="�U;mi�y
L       split_indices[$l#L       ;                                                                                                                                                                                                                    L       
split_type[$U#L       ;                                                           L       sum_hessian[$d#L       ;C��C�y�A3%CInYC	��@�TA�@CEA@��A�!B���?�i?��@��@�sB�+BӣW@�?�4@w
�@�z�AH}AB�R@M.?�/@�I?��<B�O@f�@�:bB�/�@-6?���@���?��@���A5�?���B⾋?�?�@�	?���?���B��V@�Z�?�#�@��@�\f?�w�?�1^B�Z�?�NG?��@"�?���@5��@���B���@��/L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       59L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       =:h�ʼ~�=m�;������>Y�<������>*�ǽ���=+.�>���=�r��> �����<t|>n�Ǽ�oX��==��>Q幽c�=�疽(c�>���;���<�J+�5��>�;��Nk�;�G�e�=Ps>�W<�1)�I2�.T�=��<d1�����:�>>Op���=��O��5�=�`">� ����S�?��>u���S�<�$���y>u�n;��<>)G�=�p½��ھ�1��ẍL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       =                               L       idIL       left_children[$l#L       =               	                  ��������            ��������   ����   !   #   %   '����   )   +   -����   /   1   3��������   5��������   7   9   ;��������������������������������������������������������������������������������L       loss_changes[$d#L       ==�»=�!�>vO=��>.�N;�� =��=�o�=YG�>Ŏ>/u        =�e�=��i=�OF>X?,        ><��    <�3=���>g<�=�n�    >>[%>�>a|    >i��>;'�=��h        >3��        =j��=˭�>E�                                                                                L       parents[$l#L       =���                                                           	   	   
   
                                                                                               #   #   &   &   '   '   (   (L       right_children[$l#L       =               
                  ��������            ��������    ����   "   $   &   (����   *   ,   .����   0   2   4��������   6��������   8   :   <��������������������������������������������������������������������������������L       split_conditions[$d#L       =>v�P�-��?� ?[2?�տ��@�f�W�0��g@'�?D8y=�b�<�U�=Ox�?�A�i���Iv=�=x��7�ˈ=�>�G���LD����_]=�c���o��?��=���V�`�1�@&=�<z#�=���@	bd�9$��Q2��;`�>� >?��2�`(K=x��1^�=�0����<�@)=ȍ����d�f=.���d<;7����=�uB:�|=K#3<���{m��n׻o�L       split_indices[$l#L       =                                                                                                                                                                                                                            L       
split_type[$U#L       =                                                             L       sum_hessian[$d#L       =B��;B�^�B'5PBh�$A��@-ݸBWuB\�C@EnA�0SA7`?��#?��MBwP@�#A=��B-`@��?�WAn�?���@�K@ܤAỤA�O?�(�@Am�@�Ȩ@��k?��B%�@���A��?��p?�2&@��?� @��A/T�AT�A��?��?��@!�@�;�@{�?��X?�t�B!�e?�@E�<A
�k?�@_��?��@Hq�@�p�@�@@���@"
@��tL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       61L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       #:��f���v;b/t�'�1������=��a�W"7��Qn;9�ȾSA�>���<: ?:Aߞ>�H?=��羪oW��;>$4f��~�=o���t�K=�3x�aH>���:�������>[��<a��������H��%�>m<�o{��n�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       #                  L       idIL       left_children[$l#L       #            ����   	   ��������      ����      ������������                     !��������������������������������������������L       loss_changes[$d#L       #=��y<��\=���<���    >4��>{��        >1��>-�    >Leq=ԟ4            >D�>B�>���>E�H=�9L>)�<z>                                             L       parents[$l#L       #���                                         	   	   
   
                                                      L       right_children[$l#L       #            ����   
   ��������      ����      ������������                      "��������������������������������������������L       split_conditions[$d#L       #�M��?���?�p�?sB����?���?�?�������?ڈ?A�[=�ݯ?*~V?Ώ�=�V�<�|�̅��1��>]G?� �0Y�Dl@ ��{�=��[9�����L=���;�Q��7�ν�|�=�E�;���B�L       split_indices[$l#L       #                                                                                                                              L       
split_type[$U#L       #                                   L       sum_hessian[$d#L       #C�n�@w��C��@(��?��AC���A?��?�~Y?���C��Z@E�)?���A$�C�qk?��?��@  @��@�%�C�A�=�@J��@?r@ ��@	bC{?�@�h�@���A���?�+?�X?��i?��|?�Ǣ?�)L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       35L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       !��l�:�;۽�+$�c?�>q2����h=�04:�����>��Qu�>�4��D��P��=��>&K̾�V�������%z�aY@��� >��B��=$վx�<�����b=
`? �g>�_�I��>4�i��i:L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       !                 L       idIL       left_children[$l#L       !            ����   	         ����   ��������      ������������      ����         ������������������������������������L       loss_changes[$d#L       !=��>��=�fP=�y�    >Y4>""�>��>��_    =���        >�b>���            =�3#=�S�    >�z>��=��                                    L       parents[$l#L       !���                                                     
   
                                          L       right_children[$l#L       !            ����   
         ����   ��������      ������������      ����          ������������������������������������L       split_conditions[$d#L       !?_�?T?�*F?;B=���>3�?�F�?{S����=y|?� =�?F�>���=�Qf=G�)��gͽ�͘?Q��/��Xg=�>�坾o�콕C;�k�����<1�>��=,C?�q��=Y����yL       split_indices[$l#L       !                                                                                                                           L       
split_type[$U#L       !                                 L       sum_hessian[$d#L       !C�`XC�
�A*��C�0�?�P8A��@>�C�z�@Z�p?�5V@���?�P�?�,�C�*3AJ�?�y�@��@<1@~�C�F*?�	V@���A"@7��?�*�C7�.C�%@�@��@j(�@�/�?��G?�FL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       33L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       7;���Մ<�o�.������=xw@=�Ma�м�e>X�>�� <�8>{`T�߈���<�4�C�e��C�=�b(���g>�o�=��p��Ν>�.�� =�ê>����<�s>���-�>�����=3�
<7ʾF��Y%��L>k�e=lN����=�h��D==����/�_v�-�N<*~���K>2C�<�n��6[,>�r���]L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       7                            L       idIL       left_children[$l#L       7         ����      	            ��������                  ����      !��������   #����   %����   '   )   +   -   /   1   3   5��������������������������������������������������������������������������������L       loss_changes[$d#L       7=p�
=��D=��,    =��=�V>�AN>�C=�}V>:��        =�;]:�ʀ=��M=�"=�]>3    >3�==�΀        = �G    =�L    =/�=���>W0\=���<�)�=�x=YH =�l                                                                                L       parents[$l#L       7���                                                     	   	                                                                                                     !   !   "   "L       right_children[$l#L       7         ����      
            ��������                  ����       "��������   $����   &����   (   *   ,   .   0   2   4   6��������������������������������������������������������������������������������L       split_conditions[$d#L       7��8�w����P�#����?��P� i�T�?��?� j=97 =��Z?�H�ao9�\�@UT��[P�w�ʽ����5�?z٪=��<�A��-\=!�k����<�Q3�׮�@	~���T?(Bؾ�}]�b�?]� ?�a�;[��n���'7ƽ3��=�P
<�+���<񰟼.Q�=7����9� (�P��;L�Z���=U�;ǷӽZ��=$D#���pL       split_indices[$l#L       7                                                                                                                                                                                                      L       
split_type[$U#L       7                                                       L       sum_hessian[$d#L       7B��+B63�B��d?�ԢB.l�BAibA�N�@���B��B7Ԁ@N?��NA���@�	@G�A�Z�AU�yB/�?�OVAMH\ArwN?�B?�@�@�e?�IA�I?��@s��A��B�@�)�@7�A]�@�~Al?��?�H�A]ҦA��?�>g@�@�1@6H'A�W�AY��?�N�@D�o?���?�X�?�M�A�+?њN@g_�@�&@���L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       55L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       ':u�i��ձ;a�=�3��=���>�R�:�gھ�5@�KE��|=m��=����*�
���:G�s;ux>#,>��h=�м�F;�6�=z��`��>y�������j>h�>Y�9�rOg��Y��>�_;��>nr�<�<s�>�rƾ1M>$�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       '                    L       idIL       left_children[$l#L       '            ��������   	����         ��������                           !����   #   %��������������������������������������������������������L       loss_changes[$d#L       '=���>,�>$�=rU        =�?G    =�4�><��>¸        >�>�>:6�=���=���?�z=��r=+��>a$>��    =���=Ьx                                                        L       parents[$l#L       '���                                         	   	   
   
                                                                  L       right_children[$l#L       '            ��������   
����         ��������                            "����   $   &��������������������������������������������������������L       split_conditions[$d#L       '�^��<�Ph�X �>��P=V,=���?��\��?�?}R^�/A=�G�<�RƽL��RJ\�g �=!�?�S�? I���*>��P�dR��0���?*t?�(X�@=�7N=�����bؽ�$k�:|=�؆:(�=���a��;�Y=Ɖ��n]=E�ZL       split_indices[$l#L       '                                                                                                                                          L       
split_type[$U#L       '                                       L       sum_hessian[$d#L       'C�q�@�b�C�<>@��?�O{?�eOC���@��@31^C�l�Aî�?�.U?�4f@䝟C��wA���@�SM@���@w@n�C��{Av�1?��9@�	�@>��@i.�?��?�aC?�Ū@�8?�G�?��C�y�@�AU��?��[@TF?�I�?��YL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       39L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       ��P:m����ۺU&�>V�����q=��Y:�R����k;s=��x��k>d���/�q>Y�><>��횼K����G�>X�"j�:��s�ֻy4>.�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L                    L       idIL       left_children[$l#L                   ����   	               ��������   ����������������������������   ������������L       loss_changes[$d#L       =���=�5�=�X=�e�    >Nѩ>�?=��>q�s=�GD>"r�        >�                            >'"�            L       parents[$l#L       ���                                                     	   	   
   
            L       right_children[$l#L                   ����   
               ��������   ����������������������������   ������������L       split_conditions[$d#L       ?_�?T?�*F?;B=�Ν�1�?��?7�����ƾ�rB<p�z�/N=�<�?-M�=�8W=5{~��PS�txʽ�"�=����B�?����?N�^?=Q�3L       split_indices[$l#L                                                                                                      L       
split_type[$U#L                                L       sum_hessian[$d#L       C�(wC��A$��C�&&?�ٌ@�!�@xlC��9@Pv'@��u@:hf?�?�?��AC���?ǄQ?�~p@6�?�yr@G�2?�]1?�s�C��?�,�C�Ԋ@�?�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       25L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       1; Kx�M*�<���&�Ž�+�>0<$�&�<-���;��r�>�<k�\��<� �<�	�g_K>]�����>1?3�RN>:�<e���2=�Wy��=�G\=:G�>�`L���j>��>�4.�+��1S1>��d�a�<�<B=:a��?�>��-�j��=��'>��x=�w�����: />R��>Y����L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       1                         L       idIL       left_children[$l#L       1               	            ����   ������������                  ����   !   #   %   '������������   )   +   -��������������������   /������������������������������������������������L       loss_changes[$d#L       1=R�t=�.�=��=�|>��=�vl>�'>�>T�    >e��            =�mH=��}>@%�<���>�=�cM    =~�H=�1y=���>�X            <�� =�6=���                    =ߎ!                                                L       parents[$l#L       1���                                                           
   
                                                                                 $   $L       right_children[$l#L       1               
            ����   ������������                   ����   "   $   &   (������������   *   ,   .��������������������   0������������������������������������������������L       split_conditions[$d#L       1>v�P>mf#�6��aD?�9?�zڵ�i����'\���@Ij��:�=��罄^Ⱦݑ��o��M���Nv4��_��z"�|]��X[����p���nY��ծ<ǈ�<_�K��f�����?�(=�qѺN��T�;=�k�����rC�<_H��L�=��м��L<��b=Ŵ�<����2u/�_3l=|�N=k��3twL       split_indices[$l#L       1                                                                                                                                                                                     L       
split_type[$U#L       1                                                 L       sum_hessian[$d#L       1B�
�B�Z�B#_SB���@��@��tBmdA�B�[@1@�\?�H#@��?�6!B�@��@@P�@dF�Bu�J@ ��?�Tg@3KeA���@b@�6:@O�?��?��I@��Bd�@�#�?�-�?�Å?�p?ېY?�$�A�K�?�B�?��r?�#�@ڍ?�H7?��@��BH�a?��e@W��@�~A��L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       49L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       -:��i���i;����j�>-:�ii=�c���{B�V��;� p�C+>���<�0�>;ͽ���<r�#���+=�l;���*��(:>e�5qR<
d;2L9>��؎�;:A�<�'�����j�>��v��Ϩ��6>JO��.<$�=��m�?xk=IUd�|�����<�Y��^�>ЂL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       -                       L       idIL       left_children[$l#L       -            ����   	   ����         ����   ����         ��������            !   #   %   '   )   +��������������������������������������������������������������������L       loss_changes[$d#L       -=��H=�Q�=�63=˥!    >��>J�6    =��x=��>�    >#��    =�Z/?���?P�8        >+/> -?=ނ�>�}>��>_� <� >�>M]                                                                    L       parents[$l#L       -���                                               	   	   
   
                                                                              L       right_children[$l#L       -            ����   
   ����         ����   ����         ��������             "   $   &   (   *   ,��������������������������������������������������������������������L       split_conditions[$d#L       -��n@\~?�p�N�c=5S�?���?�?����P�B��m�?A�[=��?*~V=?��|����C\��i<�N����?$��>]G>�t�?s�8��X2�ѓ�?�f����1���'2����=��[���0�5T='%��:�;E�����>9]N<q���'bq�s���n;�84���;=6-iL       split_indices[$l#L       -                                                                                                                                                                    L       
split_type[$U#L       -                                             L       sum_hessian[$d#L       -C�� AsQCC��A^�+?���C��sA*�^?�%2AJ��C�8�@@S�?��yA�/?��JA9��CDj�B�*?��7?��G@�{�@m!�@��@�˟C@�S@zK�@s�CB�q�@�)�?�H!?�z�?��N@��@=�w@J�F@O�C<Wf@�=�@3^�?��5?�S@)a�@�=B�ZN?�b�@E!�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       45L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       3������>�
rV;�E���s3i<й��/=��ҽ�A<�^v;�A��S=��!�}�B���i=�I9��P�;��J�0����>*�?=6Q��0�=��o��>`	�;��þY!F=,�<�b;�<�8���-=��˽��>i>>�����ὖL�>}>��C㺻�]�Gj>��> eN�8cμ<i���MI��K�>Z��L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       3                          L       idIL       left_children[$l#L       3               	��������               ����         ����         ����   !   #   %����   '   )   +   -   /   1��������������������������������������������������������������������������������L       loss_changes[$d#L       3=���=�@=kh�=��>0�:        >���>�3=>BW�>��=��    >�ܞ>B`>p��    >�>�p=��D    >Z�>�J=gH    >y
�=���>�>�^=�9N=�a�                                                                                L       parents[$l#L       3���                                               	   	   
   
                                                                                                L       right_children[$l#L       3               
��������               ����         ����          ����   "   $   &����   (   *   ,   .   0   2��������������������������������������������������������������������������������L       split_conditions[$d#L       3@	�F?|�G��::?*d��j���;>�-?oh>Ʉe���!??��R��c��@N�����1i��K�C��>����`��T<A?:0���M�O撽ΠԿR2�>{wݿUmj?!��[�Q���;��G�buw����=��ʉ�=�&=?�6��਼�\3=����Qw��1��oL=�X.=+�]D��bg�Ǐ���?=�*�L       split_indices[$l#L       3                                                                                                                                                                                          L       
split_type[$U#L       3                                                   L       sum_hessian[$d#L       3C��C���@.+C�\�B�T?�?�?�C��rA��1Am�A�<�C�a�?��A�#�@u��AOqP?�fAs��@��C���?���@=�A~ʷ@	~G?��A-�@���@yp�A5��@U�@T�B�(�Cm?ƨ�?�?@E|AM�?���?�g�@�h@�o@B��?��#?�h@5�Z@�m-@��?̃A?ޤ�@ɞ?���L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       51L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       ;(L�<w�l);u��>P�����=�2�<��/��n�>Z.�=[2��	P>�ͽ=4�;��M>.q
;X&���=�6N>�Y.�T�&�̙�<3Y+�d����g�;�Z>�I�(�;���=�4dL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L                       L       idIL       left_children[$l#L                      	            ����   ����   ��������   ��������������������         ����������������������������L       loss_changes[$d#L       =X�1=���=���=���=|&�=dV�=n=�m�=��"    <~�    =��R        >��                    =��>��=��Q                            L       parents[$l#L       ���                                                           
   
                              L       right_children[$l#L                      
            ����   ����   ��������   ��������������������         ����������������������������L       split_conditions[$d#L       >��^=��R?�]׻�TE>��𾾍�>�ŵ�C���]���Q�>yDb<���?���=,��cѽ�S�=QTs:��佛~�<���=��8?�1p?���?�t9̽���:.=79�I�n:�� =pL       split_indices[$l#L                                                                                                                       L       
split_type[$U#L                                      L       sum_hessian[$d#L       B�Bڐ4A@��B���@sVA�@?��B�ԇ@D?��~@��?���@���?��h?�z�B�Y�?޲�?�^?���?��^?�	]@��@i��B��u?��&@<d�?��>?˨�@�TB��B@��%L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       31L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       :X�����-;]Sƾ�d<��
>��:��=V����F�M�W=�x>Ua<��#��H�;YJ�������`�O��=�s>+î9��U�y�v�7(>��;�nо[ӥ;�>uL�9<qL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L                      L       idIL       left_children[$l#L                      	      ����   ����������������      ��������   ����      ��������������������   ��������L       loss_changes[$d#L       =��K=���=�!�=���<��<ܭ�=�\�    <D�`                =�ua>�        <{�    =忼=�U�                    >	�        L       parents[$l#L       ���                                                                                      L       right_children[$l#L                      
      ����   ����������������      ��������   ����      ��������������������   ��������L       split_conditions[$d#L       ��8\?�澣����l&>��P>`ӿi��<��a���ʼw	�= �=�	;��+?����g�D��b~���@?J�<�}�>��f�f���G�[ɬ=��G�"�����c�f�=�-�8b2�L       split_indices[$l#L                                                                                                                  L       
split_type[$U#L                                    L       sum_hessian[$d#L       C�a�@�-C��%@�3#@*�@a��C��?�ߛ@:vx?�w�?�xK?��?�Bd@�n�C��"?���?�$@BG?�-E@r��C��?�/�?�^b@��?ǭ�?�fC�l4?�x5C���L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       29L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       9��3�:��W���";��N�E��=�i���=�"X=�V'=�G� ��>"R�����g��<���:�_a���!>�]�<�iy�#l>����,�ɾ��e��"����=��M��G;�����I=��	?-e>Q0�����e�x�uV�>�>H�<W�=��ҽ�������:f<���>:ڹ�X>`E�;�hþ��a>��n��H����{=���>ͦ2=�q/�J��>�؈�C�F=�)#L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       9                             L       idIL       left_children[$l#L       9               	                  ��������         ����         !   #   %   '��������   )����   +   -��������   /   1��������   3����   5   7������������������������������������������������������������������������L       loss_changes[$d#L       9=���={��=��s>2�L>��h<��%>h{>`'�>��>�vU>X��        <~R�=���=�>�    <�1�>�G4=+W�>,MH>@8=�`0        ;���    >�2�>�        >W>�K�        ;�Հ    >Z�>�                                                                        L       parents[$l#L       9���                                                           	   	   
   
                                                                                         #   #   %   %   &   &L       right_children[$l#L       9               
                  ��������         ����          "   $   &   (��������   *����   ,   .��������   0   2��������   4����   6   8������������������������������������������������������������������������L       split_conditions[$d#L       9>]R?I��Yq`>|hv����>Pn��à>x�>���=��?��*=Bɰ�{�?��j=6��?,L��"(?@1�>�ul��de?���?Q����f���ݼ���>�����V?|?U�v=��>�ཚO">�S޻��⽓4�_%�b0?j��?%�
�,�|��߮<�&=;yӸ�%�=��(:�}���z�=�m���WE�˺�=��=��p=C�sK=�׽j�!=L       split_indices[$l#L       9                                                                                                                                                                                                            L       
split_type[$U#L       9                                                         L       sum_hessian[$d#L       9C���C�<�A*%%C�*A��@��A��C���Ab�@�AnQ�?���?���@�u�@�zC�s�?�5<@��A=��@7�'@��rA,��@�x@?��?���@��?��eC�,�@��?�4�?�"�@��&@��=?�w�?�j�@`5#?��@vW2@� I?�f�@;��?�f�?�ҿC���@�76@Li�?��@1(�?�ˆ@O��@���@�q?�d@!S�?�9@�:�?��L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       57L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       +:�y�L��<ܲ�L�/��{=�ɋ;��1�(�8=֕���MY�X���,�>g���7/�<��Z�<��d䎼��t>C�<��*=�E�=�R¾W� =8��>�����v#/>7j�;٪i�">7�]<S^��p>��˼%1�=���p�=N[��?d=���>�=�?TgL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       +                      L       idIL       left_children[$l#L       +               	               ����               ������������   ����������������������������   !   #   %��������������������   '   )������������������������L       loss_changes[$d#L       +=2փ=�=�=jm/=�)	>{=�A�=�
%=g�m=_S�    =��<�V8<���=���=���            <�S                            =�le=�y=�\                    =��Z=��                        L       parents[$l#L       +���                                                           	   	                                                         #   #   $   $L       right_children[$l#L       +               
               ����               ������������    ����������������������������   "   $   &��������������������   (   *������������������������L       split_conditions[$d#L       +���m�;*�A(��:M�5 �k� ��D�v��?��@?s����.��|a��r
�#`5��B������U��\%=j��uq<� �=�u��`�<]��=����ݽ�����B�@�>:�f=\Dp;~Q��8
z��D�=�)�?�9z@"[�S�<w���eDy<��z=��J�e�|L       split_indices[$l#L       +                                                                                                                                                          L       
split_type[$U#L       +                                           L       sum_hessian[$d#L       +B�XB���B*�uB���@ͬ�@��B��B���@g �@�U�@��@1�9@l%@CB�B��?��?�n�?��`@B�?��X?��r?� ?�3�@�)?�D�?���@mfA��nB��|?�F�?�X�?�-F?�x�?�bBA��@H�B=�A�0�A�B�A�@?�O�@�?L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       43L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       =:F���;�2��%Q=�sg����<�<����C^��U;L�N>�<�}����>b��ﯽL���J��B�����< n;?�=�Dx�rGȽ�K=^�>�Fw��Jq=}��>6-�\B	�[��=���=�"���cy<κ㽯*>T���F>+�F�Ԡ�*pX>�	=������g��}�:�XQ��q�>{� =1O>�����<oA'�� i>����f ;d#�>�9����� ��>)��L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       =                               L       idIL       left_children[$l#L       =            ����   	               ����         ����   ����         !   #   %����   '����������������   )   +   -   /   1   3   5   7   9   ;����������������������������������������������������������������������������������������L       loss_changes[$d#L       ==� O=�Uk=�=� �    >m��>�t�>��=�x>�CE>}�    >=�<�#�    <�>    >幫>E�!>E��>��>
 �    >sl                >'q�>��>/�8>e>�Q�>��>�/4?��>.�>��                                                                                        L       parents[$l#L       =���                                                     	   	   
   
                                                                                         !   !   "   "   #   #   $   $   %   %   &   &L       right_children[$l#L       =            ����   
               ����         ����   ����          "   $   &����   (����������������   *   ,   .   0   2   4   6   8   :   <����������������������������������������������������������������������������������������L       split_conditions[$d#L       =��n@�e>�	T>Ϫ�=E>>++�>�v>�?m�$����4>�=�=�-�Ⱦ|��?��|���9�ݑ����&>0��?�tN�����-�?���^E>�t�<���=�����D<�R��^<&?|)�K��Q�ξ����#v��S0��w"?�Hq>���=N4U�02Z�L��=�>J�ݲɼo��̗*9����U?=�g<#n_=�ࡽE�;��~�F�=���=4:��U=���~#���=KλL       split_indices[$l#L       =                                                                                                                                                                                                                        L       
split_type[$U#L       =                                                             L       sum_hessian[$d#L       =C��$Akx�C�D_AQ0Z?�A�CB�.B�� Ap�@z��AG��C6@c?�poB�^@�S�@	�?�~�@�b@6_yA�AC-�BB��nA+�}@)�@��G?�o?���?�C\?�9g@��t@�@+@�Y�@#��B�%C	��BlL�Ak��@��@���?�S;@E��@ �H@0�@-�@)R~@T��@
�?�g?��?B�@I'�A��B��BX.}@��C@xAKi=@�?�4J@E<�?�"L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       61L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       Y����<������.0=H|6=�&��&�{W�>��>IH�<u��>�-��ž�u=�<�=��� L->��ŽUF���r=2�T>���=+E"��%�=�N�-ܼ�|̾_r����>E�݌����>�o��qj}>���?��E�۾�:��7�> �>�ea�F�]=��5���S����W6�=�{�<'ј�a��>����<��޾G��>S�'�k���q�'��> F�=��> 
�>�@�=�kE� �L<ٍ(����=a�b����>����(���>&I�=�4�>�8>��)E>�E�=SCž`�z>�/�D%S�`�U>�l,>�%��x���"�>� U�т�?�;L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       Y                                             L       idIL       left_children[$l#L       Y               	         ����                           !   #   %   '   )   +   -   /��������   1   3   5   7   9   ;   =   ?����   A   C����   E   G   I����   K����   M��������   O   Q   S   U   W������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       Y=���>4�>��~>F�E>���>��6>���>@�-    >��?�j>���>0Z|=�$0>��>�|?���>�X>��>}�>�x�>8�x>Ȋ�>�R}>X�        >�;|>���>�>x²=� >�dP=��=�@�    =��<��n    >�Ca>�\u;��     >���    >-W�        >��>��>��h=�<L=�Q�                                                                                                                                                L       parents[$l#L       Y���                                                     	   	   
   
                                                                                                                             !   !   "   "   $   $   %   %   '   '   (   (   )   )   +   +   -   -   0   0   1   1   2   2   3   3   4   4L       right_children[$l#L       Y               
         ����                            "   $   &   (   *   ,   .   0��������   2   4   6   8   :   <   >   @����   B   D����   F   H   J����   L����   N��������   P   R   T   V   X������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       Y>w��r%@=6Z�>`Ӿچ?,��=u�ƿ��=���?M���&��h��|�=J�־4(�=���ؚ>�e��`g>�ŵ<꠼>ܙ>g����?�Z�� ľ"7?*��>
�P�&}P�T@�?��~���ܾV6=!s�Ux����������M�8����n�׾RMU���Ც�V#�� �?���?�J���=��>(�;���o��=~H��4�,�-�I�=c��=�~>�^=s��@�)<�影&c<�h���+=!��� \�:��=G��=�=�庼��=� T<}������=;��k_�����=��5=2����]�����=��f��i�fFGL       split_indices[$l#L       Y                                                                                                                                                                                                                                                                                                                             L       
split_type[$U#L       Y                                                                                         L       sum_hessian[$d#L       YC��Cbp�B�:�CB��{B5ÑB~��C>�?��AJ((Bn��A��A�<@v�Bu�vB@�&B�=A5U@��@�J�B]3�@�GAT��A0�An�?�K�?���BV�@�A�W�A���@^\_B�J(@�[{@*_?�Å@i�@`;@5�A�1�A�5B@�]?�˨A;��?�g�A�4?�-?�K�AOh(B@�@�
�@v�@�װA���@��ALH=@��?��@rA�s�B��E?�V�@���?�3?�*�?��2?��?��?���A�A�b�@+�=A��?�p�@��5@�$�@���@�8@�`AH�@�>gB2�?@W�?��{@��
?��?��@���?���L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       89L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       I;Twռ��?<�z��[�=Pi����b=v�����c�a>��y��<�;|� ��>g$<b"ս9��>S�h����au==�Ɏ��`>
�X���~�q���iu>��7=��b��D9=H)�;��ξ:��>XQ+���>F\F���2��kO<�Yk��(>S�ɽR]=B���x	{��A�=i�s���=��>�_���<=���>���l���6�>g�����;�k7����>��=ؗ���O�=��;>�9f��ތ=�!�=���ͣ>���N�<�'�3s"<M�>���=��O����L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       I                                     L       idI L       left_children[$l#L       I               	            ����                  ��������      !   #   %   '   )   +   -����   /   1   3   5��������   7��������   9����   ;   =   ?��������   A������������   C����   E   G����������������������������������������������������������������������������������������L       loss_changes[$d#L       I=h�K=��"=�5�>3F�>U�>�>\&�>+�>7��    >-1=��=���<S��=�lG>?�        >p�t=�.�>��>9:\=�O<Wsp=Hm�=<P     =u�r>5�H>&��>H�u        =�        =!'s    <�*�>=5>N�a        =+^<            =>�Z    >0��>���                                                                                        L       parents[$l#L       I���                                                           
   
                                                                                                         !   !   $   $   &   &   '   '   (   (   +   +   /   /   1   1   2   2L       right_children[$l#L       I               
            ����                  ��������       "   $   &   (   *   ,   .����   0   2   4   6��������   8��������   :����   <   >   @��������   B������������   D����   F   H����������������������������������������������������������������������������������������L       split_conditions[$d#L       I��(>�O��1���	,?ㄾmQi�QB@	�F>9��=�^�C!����>��<��>��x��F=}��򂽾q�Z��Ά�ԧҿo}�T��X�?����%[�<�v?��?�S�?#|?��p=��M����?c���Σ������Ͷ�3���g���?�r$���}���n?2h̽v<�q=�c���^<��-��fZ>q�6��]=��ɽ��N;	!���=�u.=�����v<ҷ�=��H���<��}= ]y�!Ñ=1��wK�;.�ɽWV�;*��=��_<��_���GL       split_indices[$l#L       I                                                                                                                                                                                                                                                                        L       
split_type[$U#L       I                                                                         L       sum_hessian[$d#L       IB��hB$u B���A��WA&��BK��A��A�|�@�y�@mAV�B.�[@��6@�bA��DA���?���?�y@�i@X��@�l@σ�B��@:!�@��u@Yf�?�w�@�n�A|�FA�{�@ŏm?��V?�)|@ 5?��-@8@3�?�d�@�j�A�<A���?���?�-@+��?�0`?ˈ?�E�@��i?��mAS@�W�A�'?�M�@G9�@C�5?�Q?��[?�R�?��j@3^
@%w�AL��@��UAX��@y�?���?�~�?�b`@EU�@��W@]yN@�JF@ �L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       73L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       +:_=�=��=�I��8&��D�>x�;�Zp�7�|���>f��/�/>����
{����>�M>�	Y^=����F�>}ܳ�.��.��=��;>���Bp[=�k=�y���LQ=��%>��I��4�m3�>V����@>3g��A��K��=by>�l
<�jʾ�C��n���T�`��TFL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       +                      L       idI!L       left_children[$l#L       +               	         ����               ����������������         ������������   !����   #����������������   %   '��������   )����������������������������L       loss_changes[$d#L       +=�2>��=�7A=V��=�/�>~�>^Y�='D5    >Asx=��;,) =ﴂ=Od�                <�N�<ʕ,>B��            <��.    =��j                =���>�`        =;V                             L       parents[$l#L       +���                                                     	   	   
   
                                                                 #   #L       right_children[$l#L       +               
         ����               ����������������          ������������   "����   $����������������   &   (��������   *����������������������������L       split_conditions[$d#L       +?ܭ��j��?�i��m2�g�D<G.?=�f��n�x����[���g ���?<"@=���$Ѥ<����)�?v�>�L��[�<��=̶I�iS�� L_<�^�@.`/<��=�%��r���RU�X�5�Z+z=WIG���@ ��<0ܒ=���;���Է���!ҼkA��1�L       split_indices[$l#L       +                                                                                                                                                            L       
split_type[$U#L       +                                           L       sum_hessian[$d#L       +C�8�C���AN��@^~C��@�-�@��@�?��@��C��c@.&�@L41@�ݾ?��A?���?�=`?��o@D�@C��1?��?�L
?�S_@��?�s�@���?��?��?���?�Dg@N�#C�<#?��?�G�@D�?�3�?��6?�#?�ttC���?��?��bL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       43L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       /��E1����:(�>$tU�	sX=��Z�fvȾN��<�~�>7������L����%�t�a�r<Խ�h�>�ʹ&&�>y��=�� �O�`��#(��,W>U�Q�8ƾ���F΍��4G=��>�RZ;������eSA�����T�!�W���Z
�>��<��>�>����4>���=�!>pξD�=�z'��V�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       /                        L       idI"L       left_children[$l#L       /         ����      	                     ����   ��������      ����   ������������   !   #����   %   '   )������������   +   -������������������������������������������������L       loss_changes[$d#L       /=���>u�=��    =�=f>@�>J<���=h�@>>��=�O�=�=���    <�_        =�ot=��t    =�q�            =�Sh=VU�    =$�e>=i�=��            >Kp^>^                                                L       parents[$l#L       /���                                                     	   	   
   
                                                                     !   !   "   "L       right_children[$l#L       /         ����      
                     ����   ��������      ����    ������������   "   $����   &   (   *������������   ,   .������������������������������������������������L       split_conditions[$d#L       /��#V�oͿ_�=EXg=�+�=�Kj�Vix�bd��3�r�s�C�:���`g�Tva����y+��}i=,����;�l�<���(���=�"1�D$}���V�n�w�4�þ���מ�:�9���w���[�-�ܿ0,��	��l�e�<F=�����=�ڸ<+4�=9T+�lK�=IK���;L       split_indices[$l#L       /                                                                                                                                                                        L       
split_type[$U#L       /                                               L       sum_hessian[$d#L       /C�TA,�C���?�<6@�
AA��C��b@��@'��A;�@�,a@�C�X?ɪ}@qbZ?Ƭ�?�2@�@��?�<�@:f?�R?��+?�y�C���@.I�?�1@)�@8�@�h?��?���?��@�,$C��.?�p�?�"�?�x?�Π?�0?��c@wj�?��y?���@�B)A)�C���L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       47L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       7;/��P�=Y<f����>0c�<P�F����<�h��J�<�B�<M��>����E�p<�xo=|0�	O�>��J<g����*=՛e>;�-�->3c<2i�遜>���9��=�fp��K�<�X�O'���JF=?�>k�Ծ$.I<.���>|��z<�|�=o2��{e���r��K>?8m���:�������P>����;=���؟%=��ӻv�AL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       7                            L       idI#L       left_children[$l#L       7               	                  ������������         ����      ����   !   #   %   '   )����   +��������   -   /   1������������   3������������   5��������������������������������������������������������L       loss_changes[$d#L       7=c�p=�z�=��f=���=���=�8r=�&=��>)p=�n�=��a            =��.>MR=���    >Z5�=�H0    <$h=>
!=?��=���=��f    =�;V        >eiF=�� =�!�            =uJ�            =��P                                                        L       parents[$l#L       7���                                                           	   	   
   
                                                                                         $   $   (   (L       right_children[$l#L       7               
                  ������������         ����       ����   "   $   &   (   *����   ,��������   .   0   2������������   4������������   6��������������������������������������������������������L       split_conditions[$d#L       7>v�P�-���6��W�0?�տzڵ�nTs�Iv@'�?D8y;v׮=����mH��ݑ��o��?��=��Y�=}�?���= *
>�G�?�;�X[�����p��=�щ��y
<�z�Z��&|P�ˈ?���<e9-=�SL�EX@
��:;=���>,�rC�<��̽��˼�U����=ev꺰XF��MK���=*�����<�@��=8�����L       split_indices[$l#L       7                                                                                                                                                                                                       L       
split_type[$U#L       7                                                       L       sum_hessian[$d#L       7B�d�B�d!BB\��A�{I@�LvB��A2��B/��Ah�A`�?��J@!�?�MhB%@�w@�Tz?���B)gASVO?���@��@�Ǔ@(ڨA�.�@�?�ܻ@�x@?�p�?�OB$��A��@�_�?���?�T?�L�@��i?���?�-U?��A�?�g�?��A@}��@0�@͍BM[@k!Q@��l?���@Iu<@[�n?��@�46A��
L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       55L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       +:& O�=W=�/��,�ֹv�a= Ƹ>`�.�kف<()>�B�.�> �Z�t���󻽘�a���>j]�w�<�9F>u�l�~=�P�/>� >�x�=����໺S+>OZ�;�ő�C=�]��-�Q�׼�xF>�۾ɡ����>�j�#s7�+�>߆�C[�<���L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       +                      L       idI$L       left_children[$l#L       +               	   ����   ����            ������������         ����         !��������   #   %   '   )��������������������������������������������������������L       loss_changes[$d#L       +=��=��>=l|=Ojr=�'s=�WL    ;è�    >$�A=�.�=�c�>���            <�a8>��>�C�    =�U=��=��N        > C�>�cL?#��>��O                                                        L       parents[$l#L       +���                                               	   	   
   
                                                                        L       right_children[$l#L       +               
   ����   ����            ������������         ����          "��������   $   &   (   *��������������������������������������������������������L       split_conditions[$d#L       +?ܭ��j���3�L?M$�g�D?�7=��O�m��;I���[��>��<=���-8M���G��2۽��@� �_�>�=�{A?"T�=?0��' =��5<���?��J�_o�?5�J?���4Pu=�8��j�{�ϻ��T=�e����2O�=峁�D#ܽ4[>C�jn;�hEL       split_indices[$l#L       +                                                                                                                                                             L       
split_type[$U#L       +                                           L       sum_hessian[$d#L       +C���C�6�AI��@W�C��;A5[�?�/�@��?�(;@��C�{(@���@�&-?��?�jb?�)/@At�C4�JB��@�@5A�@V:>@:?�p�?�x�@�p)C/��@ҦIB�}�?�_�?�$@G?��Z?���?�2?@J|�?�ǖ?�g3C.��@;
@j5�@�;B���L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       43L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       /���:��r����;2*�����=��~����=4j5��Bļ���(�	�Y��<�X��w;K> �����;V�a�Jvm����=�I��`+=f����>�����缯�߾�P�>�Q�cK���Խ�(��L6>R\���(T>S�Gu�=a�3>��=����2]=5���=�#��>��0=1��� ^;Va�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       /                        L       idI%L       left_children[$l#L       /               	����         ��������                  ����      ����   !   #   %   '����   )   +   -������������������������������������������������������������������������L       loss_changes[$d#L       /=��=s"9=��0=q�S<iex    =�@>)>ȕ�        <�q`=���>*�?��=��>k�)    <J}�=bN�    >$[�=�`=��P>���    >N�>ڐ>��                                                                        L       parents[$l#L       /���                                                                                                                                            L       right_children[$l#L       /               
����         ��������                  ����       ����   "   $   &   (����   *   ,   .������������������������������������������������������������������������L       split_conditions[$d#L       />]R@2xu�Yq`�`ن�T�z<����.�ӿg���_o������J�r���>���j�>��ڿ;�^�[�D�r�>��P��ƽ(sg�m�>��,#v>�*��?�0��?
X�Z���l����h�)��=|o �Kf=}7�oY�<�M�=�|�= Wy� ��<YIs�Z��D��=��<Tj��� q:��"L       split_indices[$l#L       /                                                                                                                                                                              L       
split_type[$U#L       /                                               L       sum_hessian[$d#L       /C�:C��A#�C���@1k,@��A/]A��C��~?�:y?ϛ�@�s�@g�A��>AB�9@�1�C�i�?���@J��@ȣ?��A8�@ι�@��@�N�?��(@4o;A��C��@@o�?�c?���?��@���@d,�@�u�?��@z��@*?�&<@��a?��?�n@gy�@���@���C�x�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       47L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       ';D�;�ʘ�&���,=��������0=����`�J#�>$4M=�T�+=Ey=>g�Y�f��<��:~v뾷F�>�7�;�9Q����<ƭ�=ʯҽP>� �="�<�R�) Y�_��>hcI>ދ���B=��>{*D��!�>�:�p�>�L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       '                    L       idI&L       left_children[$l#L       '      ����         	               ����         ����      ����������������      !   #��������   %��������������������������������������������L       loss_changes[$d#L       '=H�=O$�    =V�=�Y@>��>\�=�?~=��>�>b=��    >/K=���=��    =���>Y.g                =k �=���=��;        > j�                                            L       parents[$l#L       '���                                                     	   	   
   
                                                      L       right_children[$l#L       '      ����         
               ����         ����      ����������������       "   $��������   &��������������������������������������������L       split_conditions[$d#L       '?:h��K�l�.k?h�+?�V?!�T�?j�@��?J�x?��?H�=Z3�iN��fX?RX�����@IO>ѯ����E=��;�˽�+,��g�k�?��=�g<C�?��~�J�8��_#=�n�=-�ڼ�'�<>4B=������5='�F�/�=)/�L       split_indices[$l#L       '                                                                                                                                            L       
split_type[$U#L       '                                       L       sum_hessian[$d#L       'B��1B�4?��VB��B:�B��5@��A�*A�KGB~H�@{:�?�]�@�pjA�\c@&m�?�^JA��bBx�]?�ˡ@؊?���@$��@ =TA6�i@�&�?���?�@A��?��fBm+@9�?���?���A��@��@�յ?�DA'�@��L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       39L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       :4�㽰:�;X�x��c=?��>4{�:��u�q6�<��_>�an;���C�;@$��|���n�_/=�Ec�f�~;�q(�Yܕ��R
>���;v�v<�竾*����=�vL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L                     L       idI'L       left_children[$l#L                   ����   	         ������������   ����������������         ��������   ����������������L       loss_changes[$d#L       =��s=p��=�t=�Jm    =bV�=��6=��2<��            =��_                >!s>3�4=�T        =�1d                L       parents[$l#L       ���                                                                                L       right_children[$l#L                   ����   
         ������������   ����������������         ��������   ����������������L       split_conditions[$d#L       ����?ko�����>�"U<e��R~����3��z>��P=��Q;��j��Ozo�~1��L뼅�<��޿S��M��DFZ��bs=�:�>���;ܯ��L!3�׍<;.�L       split_indices[$l#L                                                                                                        L       
split_type[$U#L                                  L       sum_hessian[$d#L       C���@�MhC�ɂ@� ?��@+�	C�rf@<I/@%��?�K�?��k?���C��?�G?�KN?�?���A�̷C���Af��?��?���C�#=AF>0@�CB��B~?�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       27L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       ��s:9���N����u=٭7=o�žW9|�X����Wq>�z<�b̾3ؕ�� @>&.T=
qӾ\;�>��=S��(����}:�6ӾeO���f=����5>"� �W���EL       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L                      L       idI(L       left_children[$l#L                      	����      ����      ����      ��������������������   ����      ������������������������L       loss_changes[$d#L       =���=�oM=C$=֏�>|��    =QJ=�,�    =Z�m=��    =2�>(G�                    =��    =�i<���                        L       parents[$l#L       ���                                               	   	   
   
                              L       right_children[$l#L                      
����      ����      ����      ��������������������   ����      ������������������������L       split_conditions[$d#L       ?�2?����h�?Q�?^�<��ݿ��?p�4��
�~����;�����@?IK0=Gj�<&"1��#�=�DB<}:��н���?9��?@1½H<�O�?�@=C\���_[����L       split_indices[$l#L                                                                                                             L       
split_type[$U#L                                    L       sum_hessian[$d#L       C���C�P�@��gC��E@��`?��r@���C�!?�4�@	�a@7K`?�m@�K�C�3�?�y�?�z�?��?�M?��s@a�@5C�w@�?�z�?�ILC���@�?���?�!�L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       29L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       ;+"��6��=�`^;)�s�!Ll>plݽ�X#;�V�(�\��_�V�=�̶>�b�j��>	1.�4"<=&6:>~׽Fó<"���hђ=�ŏ�2�����>�Bֻ�i�=�Qw��7�5I�=�$L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L                       L       idI)L       left_children[$l#L                      	         ������������������������         ��������            ��������������������������������L       loss_changes[$d#L       =7�=���>G��=w')<�00<""�>N��=~1�                        =�߂=�h\=���        =��i> /=�w>#Z�                                L       parents[$l#L       ���                                                                                            L       right_children[$l#L                      
         ������������������������         ��������            ��������������������������������L       split_conditions[$d#L       ?�}�?���?5�J?:h��<�`?�_X>�I�K�l�J�	������<�(�=�C���?oM����?.G�=�g��n�q>txp�%����?��6����=+���i�{��T�=�{��B�Y��<�^kL       split_indices[$l#L                                                                                                                     L       
split_type[$U#L                                      L       sum_hessian[$d#L       B� �B״M@�ǗB�ZB@+AO@>�;@�`�B�!P?�<�?���?Ƭ�?�#�?�v�@�@��B���BŐ?��b?�DtBCjA�&A���@�eB1+2@���@���A�:eA�8A�T@a��@�9}L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       31L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       %9rY�����;)����
>=�(!>&sM: {�aJ3<�\�>�
�;�l,�{x�;t�缢U��
n���G=�1��B���L{:ȕ!=�̾��ýbr6=��L�ʅ^;l�f�].&��>�T�>-����5پ�!�=��:$��>6'�Y��>��L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       %                   L       idI*L       left_children[$l#L       %            ����   	         ��������      ����������������            ��������         !����   #������������������������������������L       loss_changes[$d#L       %=^+E=L�H=�r[=��1    =D�6=d��=GHh=!�
        =� �=��y                =�|=�H=��>�        =���>��=�d    >�[                                    L       parents[$l#L       %���                                                                                                              L       right_children[$l#L       %            ����   
         ��������      ����������������            ��������          "����   $������������������������������������L       split_conditions[$d#L       %����?�o�����>U��<����R~���n��z?^�=��b:��5�@V�@C���z ��r��^�<�~?RP<>��@ ^?*~V��(���!��~�?j�?�p佄�J�&,r=�2�=P�-��k��[�<0S9E�V=7ږ���=2�,L       split_indices[$l#L       %                                                                                                                                  L       
split_type[$U#L       %                                     L       sum_hessian[$d#L       %C���@�C�R�@���?�<:@'�?C��@B��@<�?�C?��;AM�FC���?�]z?��@?��?�@JG�A	NC�|�@�<�?��X?��n@��@���C��R?��L@)��?Ŕ�@[�A?��$?ٮ�@E&{C}R�@�{�?�??�LVL       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       37L       size_leaf_vectorSL       0}}{L       base_weights[$d#L       7����:�u���w_;����C�;Μ;�g9�EZ=̢L=_�v�:�٧�> ��+�A���;C�׾`>1>��<N��>j4>�ʽ�&z⾸�ҾR(�=��>bcý(��'4�>O�(u�>���
����|O>>׾ m>%����>��)=�P�<Ok�K�ܽ
Z��\��;���e�>r��#��I�>�"��}�>���^��=`�;�!�=��1L       
categories[$l#L        L       categories_nodes[$l#L        L       categories_segments[$L#L        L       categories_sizes[$L#L        L       default_left[$U#L       7                            L       idI+L       left_children[$l#L       7               	                           ����      ����   !   #   %   '��������������������   )����   +   -��������   /   1����   3��������   5������������������������������������������������������������L       loss_changes[$d#L       7=��=d}�=�O�>
��>ho=�=�=��>'J`>��:>|X>t$6=�=wR�>d    >��=�X    >wQ >%��;ɇ =��V                    <n�    >c�Y>�I        >bˋ>�!p    =���        =�|                                                            L       parents[$l#L       7���                                                           	   	   
   
                                                                           !   !   "   "   $   $   '   'L       right_children[$l#L       7               
                           ����       ����   "   $   &   (��������������������   *����   ,   .��������   0   2����   4��������   6������������������������������������������������������������L       split_conditions[$d#L       7>]R?I����@>|hv��>��	�>��>du�>���?��L?km?
X��ޡ�)���H=��>r�]=�R/>�9C�1�?���>��|�ݒ��|0�<�n�=��u�I�N��r=/� ��@J?�&i����,>�v�?�۲=F�&?�=���<�����b'�t�<�&���Z�:��y�=��_�D��q�h=�\���X�=�؈���<�Ɗ�((�=I�L       split_indices[$l#L       7                                                                                                                                                                                                      L       
split_type[$U#L       7                                                       L       sum_hessian[$d#L       7C��C��A�'C��\A�v�@�<�@�OTC�:.AU��A%*{A!@�G@֮@e	�?�)wC��@�f@ɵA2�d@�	@9?�@��@%j?�I�?���?��a?���@�q?���C��@���?�i�?�'@��@�ɴ?�,�@�i�?�q5?��@�A�?�8�?�y?���C��}AB�I@��?�B�@6z4@3?�@�YX?��p@hi�@ j@"7@���L       
tree_param{L       num_deletedSL       0L       num_featureSL       8L       	num_nodesSL       55L       size_leaf_vectorSL       0}}}L       nameSL       gbtree}L       learner_model_param{L       
base_scoreSL       5E-1L       boost_from_averageSL       1L       	num_classSL       3L       num_featureSL       8L       
num_targetSL       1}L       	objective{L       nameSL       multi:softprobL       softmax_multiclass_param{L       	num_classSL       3}}}L       version[#L       iii}}�2       ���R��best_iteration�Kc�best_ntree_limit�Kdubub.